`timescale 0.01 ns/1 ps
    `include "alu.v"


    module add_tb ();
        reg clock;
        reg [31:0] a, b;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] out;
        wire [49:0] pro;

        alu U1 (
                .clk(clock),
                .A(a),
                .B(b),
                .OPERATIONCODE(op),
                .O(out)
            );
        
        always
        #100 clock = ~clock; 
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clock, a, b, op, out);
            clock = 0;

    op = 3'b000;

		
		$display ("OPERATIONCODE: 000, Operation: ADD");
	
		a = 32'b10110111001001011010001101000111;
		b = 32'b01000111110110100100000110001001;
		correct = 32'b01000111110110100100000110001001;
		#400 //-9.872782e-06 * 111747.07 = 111747.07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101110110101101010101101001;
		b = 32'b01011010010101101100100000000000;
		correct = 32'b01011010010101101100100000000000;
		#400 //458927400.0 * 1.5113887e+16 = 1.5113887e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001110000100111100111101100;
		b = 32'b10011011001001011111100001111001;
		correct = 32'b11000001110000100111100111101100;
		#400 //-24.309532 * -1.3728766e-22 = -24.309532
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101111110001111000010111010;
		b = 32'b00011000000011100000110011100101;
		correct = 32'b00110101111110001111000010111010;
		#400 //1.85475e-06 * 1.835958e-24 = 1.85475e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100010110010111011101101111110;
		b = 32'b11101010101010011100110101011100;
		correct = 32'b11101010101010011100111000101000;
		#400 //-1.8790996e+21 * -1.0263912e+26 = -1.02641e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000110011000110000011101000;
		b = 32'b01010011000011001010110010000010;
		correct = 32'b01010011000011001010110010001000;
		#400 //418567.25 * 604189600000.0 = 604190000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100111000000110110010010011;
		b = 32'b10101001101111000000001000100101;
		correct = 32'b00111100111000000110110010010011;
		#400 //0.027395522 * -8.349249e-14 = 0.027395522
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011001001101101111001110100;
		b = 32'b01111011101110011100000011101010;
		correct = 32'b01111011101110011100000011101010;
		#400 //2.017322e+26 * 1.9289754e+36 = 1.9289754e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101101100111000100111010000;
		b = 32'b10100010001000001111111011100100;
		correct = 32'b00110101101100111000100111010000;
		#400 //1.3376648e-06 * -2.1818981e-18 = 1.3376648e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010101011110010010101101110011;
		b = 32'b10000110100000001001100110101001;
		correct = 32'b10010101011110010010101101110011;
		#400 //-5.0319425e-26 * -4.837403e-35 = -5.0319425e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100000011100001011000100011;
		b = 32'b10111010001101110011010001101100;
		correct = 32'b10111100000110011000100101101010;
		#400 //-0.00867227 * -0.00069887075 = -0.009371141
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110111000100001111001111101;
		b = 32'b01010001011111001010000011000100;
		correct = 32'b01010001011111001010000011000100;
		#400 //3.653151e-25 * 67814310000.0 = 67814310000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100000110101100101111100000;
		b = 32'b01110100000110111000111101111010;
		correct = 32'b01110100000110111000111101111010;
		#400 //-5.121783e-22 * 4.9299076e+31 = 4.9299076e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100010100001100011010111101;
		b = 32'b00110110101110010111000101011111;
		correct = 32'b01001100010100001100011010111101;
		#400 //54729460.0 * 5.526628e-06 = 54729460.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011100101110111101100010000;
		b = 32'b00000111000010110100110110101011;
		correct = 32'b11101011100101110111101100010000;
		#400 //-3.662579e+26 * 1.0480022e-34 = -3.662579e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010011111001010001110110110;
		b = 32'b01111101100011100111111011011000;
		correct = 32'b01111101100011100111111011011000;
		#400 //-63.159874 * 2.3676123e+37 = 2.3676123e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110000011100101011000101011;
		b = 32'b00001010011100000110011011000100;
		correct = 32'b11010110000011100101011000101011;
		#400 //-39125185000000.0 * 1.1574908e-32 = -39125185000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010110011000111011111101101;
		b = 32'b10000011001000100101000100001100;
		correct = 32'b01010010110011000111011111101101;
		#400 //439092670000.0 * -4.770056e-37 = 439092670000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010111011101010101111011101;
		b = 32'b11001011011011111011111110001010;
		correct = 32'b11101010111011101010101111011101;
		#400 //-1.4426797e+26 * -15712138.0 = -1.4426797e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110101100101000000101110111;
		b = 32'b11000010101001001011110011100111;
		correct = 32'b11111110101100101000000101110111;
		#400 //-1.186374e+38 * -82.36895 = -1.186374e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110000010000010000101011011;
		b = 32'b10001001011000100111011001000110;
		correct = 32'b11110110000010000010000101011011;
		#400 //-6.902626e+32 * -2.7259372e-33 = -6.902626e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010000011010010010100011111;
		b = 32'b00010111111101101011001101110000;
		correct = 32'b01101010000011010010010100011111;
		#400 //4.265846e+25 * 1.5942674e-24 = 4.265846e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011011111111110010010010101;
		b = 32'b11000111001001011111010001110011;
		correct = 32'b11000111001001011111010001110011;
		#400 //-3.2298225e-27 * -42484.45 = -42484.45
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011111111001001011101101101;
		b = 32'b00010010101000000000110010000000;
		correct = 32'b00011011111111001001011110010101;
		#400 //4.178776e-22 * 1.0100501e-27 = 4.178786e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011011011111000001101001001;
		b = 32'b00110010100111100101000101101001;
		correct = 32'b00110010100111100101000101101001;
		#400 //-4.6128494e-32 * 1.8430642e-08 = 1.8430642e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101111010101001100001000110;
		b = 32'b11101001011100000000011010100001;
		correct = 32'b01111101111010101001100001000110;
		#400 //3.897875e+37 * -1.8135844e+25 = 3.897875e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110111101100111001010111110111;
		b = 32'b00100111100001000110110110111001;
		correct = 32'b11110111101100111001010111110111;
		#400 //-7.2848655e+33 * 3.675632e-15 = -7.2848655e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010011101100010010010000110111;
		b = 32'b00011100101111110100111110110110;
		correct = 32'b01010011101100010010010000110111;
		#400 //1521633600000.0 * 1.2659925e-21 = 1521633600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011101101111010000100111110;
		b = 32'b00011011100000111010111111000000;
		correct = 32'b10011010110011111100010111111000;
		#400 //-3.037901e-22 * 2.1785708e-22 = -8.593303e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001111101100100001001001010;
		b = 32'b00000110001000010101100000111001;
		correct = 32'b01111001111101100100001001001010;
		#400 //1.5983119e+35 * 3.034555e-35 = 1.5983119e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011111101010010001001011000;
		b = 32'b10010010000010000101101110111010;
		correct = 32'b00011011111101010010001001000111;
		#400 //4.0554044e-22 * -4.3027095e-28 = 4.0554e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101111110010101110101000010;
		b = 32'b00101001001111001100101101110111;
		correct = 32'b00101001001111001100101101110111;
		#400 //2.3450105e-35 * 4.1920863e-14 = 4.1920863e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100011101000100010001111111;
		b = 32'b11110111000001011010100100010011;
		correct = 32'b11110111000001011010100100010011;
		#400 //0.014908909 * -2.710956e+33 = -2.710956e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000110010011111101011011000;
		b = 32'b01010010001110100011100010001101;
		correct = 32'b01010010001110100011100010001101;
		#400 //-1.4695969e-09 * 199953170000.0 = 199953170000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100011000110101001010001111;
		b = 32'b00011001011101110001101110100101;
		correct = 32'b01111100011000110101001010001111;
		#400 //4.7213035e+36 * 1.27751835e-23 = 4.7213035e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001110001101100000101100110001;
		b = 32'b10111011110001000101110100011001;
		correct = 32'b01001110001101100000101100110001;
		#400 //763546700.0 * -0.0059925434 = 763546700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001000111001111011111010101;
		b = 32'b00100110101010100101011111010010;
		correct = 32'b11011001000111001111011111010101;
		#400 //-2761412000000000.0 * 1.1819923e-15 = -2761412000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111101100101011111111101001;
		b = 32'b11001000110101100011011011010101;
		correct = 32'b11001000110101100011011011010101;
		#400 //7.570342e-20 * -438710.66 = -438710.66
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010110011010111110101100010;
		b = 32'b00010110111011000101000111100101;
		correct = 32'b10110010110011010111110101100010;
		#400 //-2.3922158e-08 * 3.817954e-25 = -2.3922158e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011111101101010101011001011;
		b = 32'b11000101100110110100000011000111;
		correct = 32'b11000101100010111101011000011010;
		#400 //493.33432 * -4968.097 = -4474.7627
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001110011010101000011101001001;
		b = 32'b00110110010111100101100101111111;
		correct = 32'b00110110010111100101100101111111;
		#400 //2.8907864e-30 * 3.3132671e-06 = 3.3132671e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010111101111000101101001001;
		b = 32'b00100000000110111001010101111100;
		correct = 32'b01110010111101111000101101001001;
		#400 //9.8062314e+30 * 1.3178471e-19 = 9.8062314e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011011100110101111101010010;
		b = 32'b10100110110111110101110100111111;
		correct = 32'b10100110110111110101110100111111;
		#400 //-7.1520704e-37 * -1.5499008e-15 = -1.5499008e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000010000000011100100010101;
		b = 32'b00110101100100010000111110011111;
		correct = 32'b11000000010000000011100100010000;
		#400 //-3.003484 * 1.0807888e-06 = -3.0034828
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001000111001001000010011100000;
		b = 32'b10100110001110111011001100111010;
		correct = 32'b10100110001110111011001100111010;
		#400 //-1.375349e-33 * -6.5121555e-16 = -6.5121555e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101000111010101100100000100;
		b = 32'b10010101111110000000110111111111;
		correct = 32'b11100101000111010101100100000100;
		#400 //-4.644085e+22 * -1.00188484e-25 = -4.644085e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000100010001110111100100011;
		b = 32'b11010010111110110001010101001110;
		correct = 32'b11110000100010001110111100100011;
		#400 //-3.3903248e+29 * -539197100000.0 = -3.3903248e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101010100000000001101001001;
		b = 32'b01001000010010010100011101001100;
		correct = 32'b01001000010010010100011101001100;
		#400 //-9.7807164e-36 * 206109.19 = 206109.19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110000000010010101001101100;
		b = 32'b11010000000001111100001010111000;
		correct = 32'b11010000000001111100001010111000;
		#400 //2.9368882e-11 * -9110741000.0 = -9110741000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011101010111000001011101100;
		b = 32'b10111111011101000101010010000101;
		correct = 32'b10111111011101000101010010000101;
		#400 //1.8595305e-17 * -0.95441467 = -0.95441467
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010011110111101011101100110;
		b = 32'b11100001101101111010100001001100;
		correct = 32'b11100001101101111010100001001100;
		#400 //3.4130874e-18 * -4.2348515e+20 = -4.2348515e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111010110010101001101000110;
		b = 32'b01011110000111100001010000010001;
		correct = 32'b01011111100000000110110000100101;
		#400 //1.5659937e+19 * 2.847687e+18 = 1.8507624e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000111100000010100010001111;
		b = 32'b10111011101001001011110101001100;
		correct = 32'b10111011101001001011110101001100;
		#400 //1.445401e-33 * -0.0050274488 = -0.0050274488
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101010110111110011111000011;
		b = 32'b01101100001101001011111010111011;
		correct = 32'b01101100001101001011101101001011;
		#400 //-6.4904594e+22 * 8.740294e+26 = 8.7396445e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111100110000110011100100111;
		b = 32'b11011011110101011100110111000011;
		correct = 32'b11011011110101011100110111000011;
		#400 //1.8167846e-05 * -1.20360815e+17 = -1.20360815e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100100010111100000001101011;
		b = 32'b11100110110111101111110011001100;
		correct = 32'b01110100100010111100000001101011;
		#400 //8.857812e+31 * -5.2651432e+23 = 8.857812e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001001100111111110100101000;
		b = 32'b00010000000000001001100101001011;
		correct = 32'b11111001001100111111110100101000;
		#400 //-5.8409735e+34 * 2.5361642e-29 = -5.8409735e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000110011111101101010000100;
		b = 32'b01101110111010011011100011100000;
		correct = 32'b11110000110000010011111011110110;
		#400 //-5.1462053e+29 * 3.6166754e+28 = -4.7845378e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011000101011011011001100111;
		b = 32'b11011010011001101000011000011011;
		correct = 32'b11111011000101011011011001100111;
		#400 //-7.773518e+35 * -1.6221674e+16 = -7.773518e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001100001100110010101001010;
		b = 32'b01011000011110010111011001100101;
		correct = 32'b01011000011110010111001000110010;
		#400 //-72153120000.0 * 1097147600000000.0 = 1097075440000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011000011001100100011000100;
		b = 32'b00111100011001111000011011001000;
		correct = 32'b01011011000011001100100011000100;
		#400 //3.962724e+16 * 0.014131255 = 3.962724e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100001100011110101100000111;
		b = 32'b00001101011110100001111101001110;
		correct = 32'b10111100001100011110101100000111;
		#400 //-0.010859258 * 7.707488e-31 = -0.010859258
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011110101010110100001101010;
		b = 32'b10100011110110111111110111000011;
		correct = 32'b00111011110101010110100001101010;
		#400 //0.0065126913 * -2.38515e-17 = 0.0065126913
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111100001011111100010110010;
		b = 32'b11001010101101000101001101100101;
		correct = 32'b11001010101101000101001101100101;
		#400 //3.718455e-15 * -5908914.5 = -5908914.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000101001111110011101111110;
		b = 32'b11010001100010100001000110101010;
		correct = 32'b11010001100010100001000110000000;
		#400 //343867.94 * -74125230000.0 = -74124890000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000011010110011000101101110;
		b = 32'b10000101101101101111011100111100;
		correct = 32'b00110000011010110011000101101110;
		#400 //8.5562746e-10 * -1.7206017e-35 = 8.5562746e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000000101011000100010000001;
		b = 32'b11100101100101010110111011111111;
		correct = 32'b11100101100101010110111011111111;
		#400 //-153122.02 * -8.8210015e+22 = -8.8210015e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011000110010111010010110111;
		b = 32'b10011010011010011100010000111101;
		correct = 32'b11100011000110010111010010110111;
		#400 //-2.830762e+21 * -4.834179e-23 = -2.830762e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010000000101110100101110000;
		b = 32'b01011100110010111011000011100001;
		correct = 32'b01011100110010111011000011100001;
		#400 //9.617885e-38 * 4.586712e+17 = 4.586712e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110000100111110001111101110;
		b = 32'b00000000110000001011111100111111;
		correct = 32'b01101110000100111110001111101110;
		#400 //1.1442462e+28 * 1.7701021e-38 = 1.1442462e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100110100000101011001111111;
		b = 32'b11010100010000010000101101001011;
		correct = 32'b01100100110100000101011001111111;
		#400 //3.0745244e+22 * -3316472600000.0 = 3.0745244e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000111101110111011110000100;
		b = 32'b10000101110011000001101110000110;
		correct = 32'b11010000111101110111011110000100;
		#400 //-33214440000.0 * -1.9194178e-35 = -33214440000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111001101011100011000001100;
		b = 32'b01000101101111111000111010010110;
		correct = 32'b01100111001101011100011000001100;
		#400 //8.5840165e+23 * 6129.823 = 8.5840165e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111111100101000000000001110;
		b = 32'b00100001001000110011011011110100;
		correct = 32'b00100001001000110011011100010010;
		#400 //1.5671209e-24 * 5.529928e-19 = 5.5299433e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101010111010011111110010000;
		b = 32'b11001100100010101110110010110101;
		correct = 32'b11001100100010101110110010110101;
		#400 //0.054015696 * -72836520.0 = -72836520.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110101011011011010111000010;
		b = 32'b00111001100011011101111010011101;
		correct = 32'b00111001100011011101111010011010;
		#400 //-7.899416e-11 * 0.00027059476 = 0.00027059467
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001101000100001001010001110;
		b = 32'b01010001000101000111011001111010;
		correct = 32'b01010001000101000111011001111010;
		#400 //3.901753e-33 * 39852680000.0 = 39852680000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111000111100001100000000000;
		b = 32'b10010111011001111111010101100000;
		correct = 32'b10100111000111100001100000000000;
		#400 //-2.1939915e-15 * -7.494983e-25 = -2.1939915e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010001000101100011111011100;
		b = 32'b11000101000101101110010011010000;
		correct = 32'b11000101000101101110010011010000;
		#400 //-5.136453e-28 * -2414.3008 = -2414.3008
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010011011111111110100100011;
		b = 32'b11001101010010010101001101001110;
		correct = 32'b11001101010010010101001101010010;
		#400 //-59.997204 * -211105000.0 = -211105060.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110100000110111101011001010;
		b = 32'b11001110111100011100010101100100;
		correct = 32'b11001110111100011100010011100001;
		#400 //16829.395 * -2028122600.0 = -2028105900.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000111100011001101011111010;
		b = 32'b10001010011010111101011011100110;
		correct = 32'b11011000111100011001101011111010;
		#400 //-2125183400000000.0 * -1.1355256e-32 = -2125183400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101010000010011011100110100101;
		b = 32'b00001110010101000010000101111101;
		correct = 32'b00101010000010011011100110100101;
		#400 //1.2232453e-13 * 2.6147142e-30 = 1.2232453e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110000101101110110001110110;
		b = 32'b00100011110110010110001100010011;
		correct = 32'b00100011110110010110001100010011;
		#400 //2.8385588e-35 * 2.3569147e-17 = 2.3569147e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110010010111000110101011110;
		b = 32'b00001001111000001000000010000001;
		correct = 32'b01011110010010111000110101011110;
		#400 //3.6668707e+18 * 5.4046883e-33 = 3.6668707e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011111111110100011111000110;
		b = 32'b10011111110101110010110001101100;
		correct = 32'b01100011111111110100011111000110;
		#400 //9.418183e+21 * -9.112953e-20 = 9.418183e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101100100000000000000101011;
		b = 32'b01100000011011000001010111101000;
		correct = 32'b01100000011011000001010111101000;
		#400 //2.4980132e-16 * 6.8047033e+19 = 6.8047033e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010001000000010000001100000;
		b = 32'b10100000000010000110101110011001;
		correct = 32'b11101010001000000010000001100000;
		#400 //-4.8395254e+25 * -1.1555249e-19 = -4.8395254e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101110100001111110010000111;
		b = 32'b01011010001111100110010110001110;
		correct = 32'b01110101110100001111110010000111;
		#400 //5.2984356e+32 * 1.3397977e+16 = 5.2984356e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000111010111100101111111111110;
		b = 32'b01010010111110110011011001101100;
		correct = 32'b01010010111110110011011001101100;
		#400 //-1.6729633e-34 * 539474920000.0 = 539474920000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111001100101001011100011000;
		b = 32'b11010000111110010000101001010011;
		correct = 32'b11010000111110010000101001010011;
		#400 //3.7817948e-20 * -33425627000.0 = -33425627000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111110000010110110110011010;
		b = 32'b10101000100010111010111000011111;
		correct = 32'b10101000100010111010111000011111;
		#400 //2.910383e-34 * -1.5507613e-14 = -1.5507613e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010001101110010000111000001;
		b = 32'b10000001100000010101011111010011;
		correct = 32'b10110010001101110010000111000001;
		#400 //-1.0659677e-08 * -4.751314e-38 = -1.0659677e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100011100000100101001011011;
		b = 32'b11011010110111111100101110100110;
		correct = 32'b01110100011100000100101001011011;
		#400 //7.6151084e+31 * -3.1496417e+16 = 7.6151084e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101000010010000000111101110;
		b = 32'b00100101010011011100011110100101;
		correct = 32'b01110101000010010000000111101110;
		#400 //1.7367769e+32 * 1.7848558e-16 = 1.7367769e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111000010001111111110111110;
		b = 32'b11001011100100000100010010100101;
		correct = 32'b11001011100100000100010010100101;
		#400 //-6.754572e-30 * -18909514.0 = -18909514.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100100000001100000101100001;
		b = 32'b11111111001111001001100111110010;
		correct = 32'b11111111001110001001001111100111;
		#400 //5.3482895e+36 * -2.506942e+38 = -2.453459e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010011110010111100011011011;
		b = 32'b11100010010110010110011101010110;
		correct = 32'b11100010010110010110011101010110;
		#400 //-1.4521187e-08 * -1.0025974e+21 = -1.0025974e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100100101001101101100110010;
		b = 32'b00101011011101100001111100111011;
		correct = 32'b00101011011101100001111100111011;
		#400 //2.2934934e-31 * 8.74401e-13 = 8.74401e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111010011000101110101000000010;
		b = 32'b01000110110001100110110101110100;
		correct = 32'b11111010011000101110101000000010;
		#400 //-2.9455133e+35 * 25398.727 = -2.9455133e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010010011011101110000010100;
		b = 32'b00011010110110111001111001000001;
		correct = 32'b10111010010011011101110000010100;
		#400 //-0.00078529236 * 9.083195e-23 = -0.00078529236
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100110000010101110100110011;
		b = 32'b11000011011001110011100000010010;
		correct = 32'b11000011011001110011100000010010;
		#400 //-1.952478e-26 * -231.21902 = -231.21902
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110100110100101001000110010;
		b = 32'b11110110110100101110001011010000;
		correct = 32'b11110110110100101110001011010000;
		#400 //5.8049137e-35 * -2.138638e+33 = -2.138638e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010000101000001000111011001;
		b = 32'b10010010001111101111010101011000;
		correct = 32'b00100010000101000001000111011001;
		#400 //2.0067189e-18 * -6.025584e-28 = 2.0067189e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110000111111000111111010101;
		b = 32'b01110110010100001111010011011010;
		correct = 32'b01110110010100001111010011011010;
		#400 //-1.2889303e-25 * 1.0595351e+33 = 1.0595351e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100010010101001111001001101;
		b = 32'b00001010010000001100010010101000;
		correct = 32'b11000100010010101001111001001101;
		#400 //-810.47345 * 9.281451e-33 = -810.47345
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101000011000110000100111111;
		b = 32'b00111101101011001001100011001101;
		correct = 32'b11111101000011000110000100111111;
		#400 //-1.1662303e+37 * 0.08427582 = -1.1662303e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100010000111010010000000100111;
		b = 32'b11110100110010111000101100101011;
		correct = 32'b11110100110010111000101100101011;
		#400 //-7.246139e+20 * -1.290111e+32 = -1.290111e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011111110100100110111100111;
		b = 32'b00001000000010100011110101111000;
		correct = 32'b11101011111110100100110111100111;
		#400 //-6.0519868e+26 * 4.160012e-34 = -6.0519868e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001011000100101110000100111;
		b = 32'b00101010100101100001001111010101;
		correct = 32'b01100001011000100101110000100111;
		#400 //2.6097528e+20 * 2.6659114e-13 = 2.6097528e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111010000010111110100111011;
		b = 32'b00010010011001010010111000110111;
		correct = 32'b11000111010000010111110100111011;
		#400 //-49533.23 * 7.2316623e-28 = -49533.23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000111000011011101100110111;
		b = 32'b00011110000110100101000010111011;
		correct = 32'b00011110000110100011010010000100;
		#400 //-5.8350176e-24 * 8.169387e-21 = 8.163552e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111001000011001110001100111;
		b = 32'b01001000100111000110110100100111;
		correct = 32'b11001111001000011001011110000100;
		#400 //-2711381800.0 * 320361.22 = -2711061500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010011001010101001111111011;
		b = 32'b00100100101011011111110111110110;
		correct = 32'b10111010011001010101001111111011;
		#400 //-0.0008748171 * 7.545702e-17 = -0.0008748171
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000011111011001011111110011100;
		b = 32'b11100101111100010011000110110001;
		correct = 32'b11100101111100010011000110110001;
		#400 //-473.49695 * -1.4237587e+23 = -1.4237587e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010100010010010011010010001;
		b = 32'b10010110101001010101001110111100;
		correct = 32'b01101010100010010010011010010001;
		#400 //8.290248e+25 * -2.6710032e-25 = 8.290248e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101101100010110111010101010;
		b = 32'b01101010100001100000101000110000;
		correct = 32'b01101101101100111000011011010011;
		#400 //6.864079e+27 * 8.102208e+25 = 6.945101e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101101100111011110011011111;
		b = 32'b01011100010010100001101010100000;
		correct = 32'b01110101101100111011110011011111;
		#400 //4.556894e+32 * 2.2754888e+17 = 4.556894e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000011101000000111101010010;
		b = 32'b00010101001111011011101101010010;
		correct = 32'b10110000011101000000111101010010;
		#400 //-8.8788454e-10 * 3.8316016e-26 = -8.8788454e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101100010110011101010100110;
		b = 32'b11111111011001101110111011111010;
		correct = 32'b11111111011001101110111011111010;
		#400 //-2.4152398e-16 * -3.0696328e+38 = -3.0696328e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100000101111111101111111100;
		b = 32'b00111101000100010001111111001011;
		correct = 32'b11111100000101111111101111111100;
		#400 //-3.1565907e+36 * 0.03543071 = -3.1565907e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101100111111111010001011011;
		b = 32'b00011010010001011011100101110110;
		correct = 32'b00111101100111111111010001011011;
		#400 //0.07810279 * 4.088846e-23 = 0.07810279
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010000001011011011111011110;
		b = 32'b11001110110010101111001111001101;
		correct = 32'b01011010000001011011011111011100;
		#400 //9409584000000000.0 * -1702487700.0 = 9409582000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011100111101110111110010001111;
		b = 32'b10110000111110110101000011101110;
		correct = 32'b10110000111110110101000011101110;
		#400 //1.6377287e-21 * -1.8285655e-09 = -1.8285655e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001111000010000010110100110;
		b = 32'b01110111111110000000101011010101;
		correct = 32'b01110111111110000000101011010101;
		#400 //-3.5502222e-28 * 1.00617916e+34 = 1.00617916e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100111001000000011011101110;
		b = 32'b10111110010010010111101110101000;
		correct = 32'b11011100111001000000011011101110;
		#400 //-5.134713e+17 * -0.19676077 = -5.134713e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111111101101000001011111100;
		b = 32'b10011100110011010001011100010011;
		correct = 32'b01001111111101101000001011111100;
		#400 //8271558700.0 * -1.3571727e-21 = 8271558700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001100011000111111110111100;
		b = 32'b00101100100011110000000010000100;
		correct = 32'b11011001100011000111111110111100;
		#400 //-4943368000000000.0 * 4.0643617e-12 = -4943368000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001000011001111011001001010;
		b = 32'b01101100100100111110001001111100;
		correct = 32'b01101100100100111110001001111100;
		#400 //-2.051268e-09 * 1.4302531e+27 = 1.4302531e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110101010011010000111111111001;
		b = 32'b10100110001110111010011010010110;
		correct = 32'b11110101010011010000111111111001;
		#400 //-2.5994747e+32 * -6.5104424e-16 = -2.5994747e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110001000011111110010000010;
		b = 32'b00011000001110100100101101000110;
		correct = 32'b11000110001000011111110010000010;
		#400 //-10367.127 * 2.407794e-24 = -10367.127
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000000000111101111000110011;
		b = 32'b00101100111001010010001111111111;
		correct = 32'b01110000000000111101111000110011;
		#400 //1.6324463e+29 * 6.512568e-12 = 1.6324463e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100110111001101101100010001;
		b = 32'b00010010001011111101111001001110;
		correct = 32'b10111100110111001101101100010001;
		#400 //-0.026959928 * 5.5494275e-28 = -0.026959928
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001001101110010101111011100;
		b = 32'b10011110011101101110001001111010;
		correct = 32'b10011110011101101110001001111010;
		#400 //-3.364326e-38 * -1.3069966e-20 = -1.3069966e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011101110000011111111001101;
		b = 32'b01110001000100111101001011010000;
		correct = 32'b01110001000100111101001011010000;
		#400 //3.0481477e-22 * 7.3198645e+29 = 7.3198645e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010011100000010010110100000;
		b = 32'b00110111001100010011000010100100;
		correct = 32'b11011010011100000010010110100000;
		#400 //-1.6898841e+16 * 1.0561347e-05 = -1.6898841e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011101011000100011011110101;
		b = 32'b01100001011010100100001010011111;
		correct = 32'b01100001011010100100001010011111;
		#400 //1.224103e-12 * 2.7008367e+20 = 2.7008367e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001001001001100001001111100;
		b = 32'b10101101111000110110011000111111;
		correct = 32'b01001001001001001100001001111100;
		#400 //674855.75 * -2.5852319e-11 = 674855.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101001011111100110111100110;
		b = 32'b11000011011001100100110011001000;
		correct = 32'b11010101001011111100110111100110;
		#400 //-12081179000000.0 * -230.29993 = -12081179000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010110000110101111101111000;
		b = 32'b01101000010000101111101110110100;
		correct = 32'b01101000010000101111101110110100;
		#400 //-5.2955937e-18 * 3.6831288e+24 = 3.6831288e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010000111001000110000100010;
		b = 32'b00010111111101100001011011001011;
		correct = 32'b01110010000111001000110000100010;
		#400 //3.1007406e+30 * 1.5903131e-24 = 3.1007406e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111111010000000110001110111;
		b = 32'b01111011111000001101010011111001;
		correct = 32'b01111011111000001101010011111001;
		#400 //1.8128804 * 2.3347882e+36 = 2.3347882e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100100000100111010011011001;
		b = 32'b01110001011111101010110000100100;
		correct = 32'b01110001011111101010110000100100;
		#400 //-1043.6515 * 1.2610768e+30 = 1.2610768e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110010101000110000111000000;
		b = 32'b11001100111101101110011000001100;
		correct = 32'b11010110010101000110000111011111;
		#400 //-58379075000000.0 * -129445980.0 = -58379205000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110110101111001001011100000;
		b = 32'b10011110101011111111100111000100;
		correct = 32'b10111110110101111001001011100000;
		#400 //-0.42104244 * -1.8632146e-20 = -0.42104244
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001011011101101000111101100;
		b = 32'b11000110111000010010001000001110;
		correct = 32'b11000110111000010010001000001110;
		#400 //-3.4752885e-09 * -28817.027 = -28817.027
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101100100010010110001001000;
		b = 32'b00000011110001011001011001100000;
		correct = 32'b00110101100100010010110001001000;
		#400 //1.0816229e-06 * 1.1613144e-36 = 1.0816229e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011011101010010010101001110;
		b = 32'b01000000000101010000001000001101;
		correct = 32'b01001011011101010010010101010000;
		#400 //16065870.0 * 2.3282502 = 16065872.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110011001011000000001000111;
		b = 32'b00000001000100010001110111110101;
		correct = 32'b11011110011001011000000001000111;
		#400 //-4.134324e+18 * 2.6653787e-38 = -4.134324e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111001101001001100111111111;
		b = 32'b01011011000110111101111010110111;
		correct = 32'b01011011000110111101111010110111;
		#400 //-8.904344e-30 * 4.38735e+16 = 4.38735e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101100011011011111000100110;
		b = 32'b00011110101010010100100000110110;
		correct = 32'b00100101100011011100000011001011;
		#400 //2.458845e-16 * 1.7923437e-20 = 2.4590243e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010001010000001110101111100;
		b = 32'b11001010001111111011100001011111;
		correct = 32'b11011010001010000001110101111100;
		#400 //-1.1830054e+16 * -3141143.8 = -1.1830054e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111111001010101101110110000;
		b = 32'b00100111101111010000000111110111;
		correct = 32'b10111111111001010101101110110000;
		#400 //-1.7918606 * 5.246017e-15 = -1.7918606
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001100111110000110110101111;
		b = 32'b00110011110101010111000111010001;
		correct = 32'b11001001100111110000110110101111;
		#400 //-1302965.9 * 9.9392885e-08 = -1302965.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100000000001101101001100011;
		b = 32'b01001110110110111010101011111000;
		correct = 32'b01001110110110111010101011111000;
		#400 //-4.2633906e-22 * 1842707500.0 = 1842707500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101001011101111100000000011;
		b = 32'b01101100011111010001011111110000;
		correct = 32'b01101100011111010001011111110000;
		#400 //8.226993e-36 * 1.2238851e+27 = 1.2238851e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010100101111001100001111110111;
		b = 32'b01111101101001011010010001001011;
		correct = 32'b01111101101001011010010001001011;
		#400 //1.9060443e-26 * 2.752196e+37 = 2.752196e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101110011000011011111101100;
		b = 32'b10101000001000010010000111101000;
		correct = 32'b10101101110011000100110000010000;
		#400 //-2.321695e-11 * -8.944648e-15 = -2.3225893e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001101010111001111001001110;
		b = 32'b10110101010101111001100011101010;
		correct = 32'b10110101010101111001100011101001;
		#400 //7.621387e-14 * -8.031626e-07 = -8.0316255e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111110101000011101011110000;
		b = 32'b01111001100111111110011000101010;
		correct = 32'b01111001100111111110011000101010;
		#400 //-2.0044578e+24 * 1.0378044e+35 = 1.0378044e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000010000110111010000000000010;
		b = 32'b01110110000100000100100111010100;
		correct = 32'b01110110000100000100100111010100;
		#400 //-1.1433522e-37 * 7.316291e+32 = 7.316291e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010110101101010111001111101;
		b = 32'b01110011110100111111100000000010;
		correct = 32'b01110011110100111111100000000010;
		#400 //3.1544625e-37 * 3.3587794e+31 = 3.3587794e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000111011010011100001110011;
		b = 32'b10110000111111010001000001110000;
		correct = 32'b10110000111111010001000001110000;
		#400 //-6.1320063e-24 * -1.8412845e-09 = -1.8412845e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101110111100100010000100111;
		b = 32'b11101000100001010101011000110000;
		correct = 32'b11101000100001010101011000110000;
		#400 //-1.6560124e-06 * -5.037317e+24 = -5.037317e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100010001101110000010000110;
		b = 32'b01001110011110000100101011100001;
		correct = 32'b01001110011110000100101011100001;
		#400 //-6.5802894e-22 * 1041414200.0 = 1041414200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110011110100001110111111010;
		b = 32'b10010111101001011110101111010010;
		correct = 32'b00110110011110100001110111111010;
		#400 //3.7270352e-06 * -1.07224045e-24 = 3.7270352e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101100111001010000101010100;
		b = 32'b01000110111100110100000000010111;
		correct = 32'b01011101100111001010000101010100;
		#400 //1.4107993e+18 * 31136.045 = 1.4107993e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010010100101110010001100000;
		b = 32'b11001010011010000001111100100100;
		correct = 32'b11001010011010000001111100100100;
		#400 //4.3611462e-23 * -3803081.0 = -3803081.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111000110101111111010100001001;
		b = 32'b00110011101100010001000100100011;
		correct = 32'b01111000110101111111010100001001;
		#400 //3.5041054e+34 * 8.245322e-08 = 3.5041054e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011011110000110111111111101;
		b = 32'b11010100011111000111001110000101;
		correct = 32'b11010100011111000111001110000101;
		#400 //5.7843852e-08 * -4337079400000.0 = -4337079400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000011011101110101001000100100;
		b = 32'b10110001100100111110010101000010;
		correct = 32'b10110001100100111110010101000010;
		#400 //7.268107e-37 * -4.3043267e-09 = -4.3043267e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101111110001100100111001011;
		b = 32'b00110001000100111101101110001101;
		correct = 32'b11101101111110001100100111001011;
		#400 //-9.6245294e+27 * 2.1516116e-09 = -9.6245294e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101001010101110010110011110;
		b = 32'b11000001000011011111001111000001;
		correct = 32'b11000001000011011111001111000001;
		#400 //-8.0355356e-36 * -8.87201 = -8.87201
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110111010100011011010110000;
		b = 32'b11101101111111011011001110110111;
		correct = 32'b11101101111111011011001110110111;
		#400 //8.438435e+18 * -9.814621e+27 = -9.814621e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110100101111000001110011001;
		b = 32'b01100001000001000010101011010110;
		correct = 32'b01100001000001000010101011010110;
		#400 //-2.4478416e-25 * 1.5237855e+20 = 1.5237855e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100101010100101101000101001;
		b = 32'b01101101000011101001111101011000;
		correct = 32'b01101101000011101001111101011000;
		#400 //-5853256600000.0 * 2.758719e+27 = 2.758719e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001100100000111111100000101;
		b = 32'b11011110000101111011110001000100;
		correct = 32'b11100001100100011010111001111110;
		#400 //-3.331855e+20 * -2.7334222e+18 = -3.3591892e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101100101000011011011011110111;
		b = 32'b11011010000111011110011101011011;
		correct = 32'b11011010000111011110011101011011;
		#400 //-4.5962084e-12 * -1.1111487e+16 = -1.1111487e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011101001111011111111111000;
		b = 32'b01111110000010010000101100000001;
		correct = 32'b01111110000010010000101100000001;
		#400 //-2.775189e-22 * 4.5540343e+37 = 4.5540343e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000100011100110001000101111110;
		b = 32'b11110101111000101001100011110010;
		correct = 32'b11110101111000101001100011110010;
		#400 //2.8572545e-36 * -5.7449277e+32 = -5.7449277e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101111000111010110011100000;
		b = 32'b11110001010011011110011000110001;
		correct = 32'b11110001010011011110011000101111;
		#400 //1.3439577e+23 * -1.0195634e+30 = -1.0195632e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001100011011001000110101011;
		b = 32'b01011101100111000001100100100010;
		correct = 32'b01011101100111000001100100100010;
		#400 //2.2335652e-28 * 1.4060074e+18 = 1.4060074e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110101100100011001010100010;
		b = 32'b00011100100001101011111100100100;
		correct = 32'b11001110101100100011001010100010;
		#400 //-1494831400.0 * 8.916785e-22 = -1494831400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011001011101111101001010000;
		b = 32'b11000110000000010000111010000011;
		correct = 32'b11001011001011110001101010010100;
		#400 //-11467344.0 * -8259.628 = -11475604.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110001010010110000011010111;
		b = 32'b01011001011110001110110110100101;
		correct = 32'b01011001011110001110110110100101;
		#400 //2.523933e-06 * 4379193000000000.0 = 4379193000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000000110011011111000011100;
		b = 32'b11101001011000101111101110000010;
		correct = 32'b01110000000110011011101010010000;
		#400 //1.9032414e+29 * -1.7150309e+25 = 1.9030699e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010010000011101011110011110;
		b = 32'b10101011000001111000101101110010;
		correct = 32'b11101010010000011101011110011110;
		#400 //-5.8585227e+25 * -4.8155154e-13 = -5.8585227e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110010101000100111110110100;
		b = 32'b11111100000001110000111100101111;
		correct = 32'b11111100000001110000111100101111;
		#400 //-13587.926 * -2.805072e+36 = -2.805072e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100101001000000110001101111;
		b = 32'b00100100011111101010010010011010;
		correct = 32'b01100100101001000000110001101111;
		#400 //2.4209296e+22 * 5.5216893e-17 = 2.4209296e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001111000111110101111001000;
		b = 32'b00000100110000101101101100111011;
		correct = 32'b11011001111000111110101111001000;
		#400 //-8019258000000000.0 * 4.5810512e-36 = -8019258000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110101010100100101100001100;
		b = 32'b01001001101100010001100011000010;
		correct = 32'b01001001101100111100000111101110;
		#400 //21797.523 * 1450776.2 = 1472573.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001100001101100110110111100;
		b = 32'b01111111010000101010010000111011;
		correct = 32'b01111111010000101010010000111011;
		#400 //-4.951904e-38 * 2.5872296e+38 = 2.5872296e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010110110111000110010001001;
		b = 32'b10100010011111100100000110110100;
		correct = 32'b00110010110110111000110010001001;
		#400 //2.5558863e-08 * -3.4458202e-18 = 2.5558863e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000001101001111011110111011;
		b = 32'b10001101001100101101110011011101;
		correct = 32'b01010000001101001111011110111011;
		#400 //12144537000.0 * -5.511634e-31 = 12144537000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000111001110111100111111101;
		b = 32'b10001100001000011111011010001101;
		correct = 32'b10100000111001110111100111111101;
		#400 //-3.9213647e-19 * -1.2477183e-31 = -3.9213647e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110110111010101010001110100;
		b = 32'b00110110011001111110100001111010;
		correct = 32'b00111110110111010101010011101000;
		#400 //0.43228495 * 3.4557002e-06 = 0.4322884
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111000110001000000101010110;
		b = 32'b01001001100011000000001101001111;
		correct = 32'b01001001100100001100011101011010;
		#400 //39041.336 * 1146985.9 = 1186027.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000110101001000100001110010100;
		b = 32'b10111100100111010101011011101011;
		correct = 32'b10111100100111010101011011101011;
		#400 //-6.178924e-35 * -0.019206485 = -0.019206485
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110101000001000100111110001;
		b = 32'b01110101110000000000100110001001;
		correct = 32'b01110101110000000000100110001001;
		#400 //2.5936447e-25 * 4.8687226e+32 = 4.8687226e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001111100110100001101001000;
		b = 32'b11000010000011100000100001001011;
		correct = 32'b11000010100000111101010011111000;
		#400 //-30.407852 * -35.5081 = -65.915955
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111001000110111111001101110110;
		b = 32'b00011100010111110011101100000110;
		correct = 32'b10111001000110111111001101110110;
		#400 //-0.00014872648 * 7.3860797e-22 = -0.00014872648
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010111011001000100110010111;
		b = 32'b01101001100111100111000011111000;
		correct = 32'b01101001100111100111000011111000;
		#400 //507960330000.0 * 2.394297e+25 = 2.394297e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110111001000101111110010000;
		b = 32'b10110100100111010100111011110100;
		correct = 32'b11110110111001000101111110010000;
		#400 //-2.3159803e+33 * -2.9300975e-07 = -2.3159803e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100001000010101000000110101110;
		b = 32'b01010011000010101000111010101101;
		correct = 32'b01010011000010101000111010101101;
		#400 //-4.692785e-19 * 595099200000.0 = 595099200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110001001111000010011010010100;
		b = 32'b11011001100011011001100110011010;
		correct = 32'b01110001001111000010011010010100;
		#400 //9.316771e+29 * -4982107300000000.0 = 9.316771e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110010111100000001000000001;
		b = 32'b01000101011000000011111011000000;
		correct = 32'b01000101011000000011111011000000;
		#400 //5.0478736e-11 * 3587.9219 = 3587.9219
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101100001101101111100111111;
		b = 32'b00010001011000101110110100001011;
		correct = 32'b01000101100001101101111100111111;
		#400 //4315.906 * 1.7901301e-28 = 4315.906
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001101001000101111111001011;
		b = 32'b11101110011010010101001111001011;
		correct = 32'b11101110011010010101001111001011;
		#400 //4.7839186e-09 * -1.8052827e+28 = -1.8052827e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001111010100010111001111001;
		b = 32'b10011000001100110011011100010000;
		correct = 32'b01001001111010100010111001111001;
		#400 //1918415.1 * -2.3163007e-24 = 1918415.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010010011011000000000000000;
		b = 32'b11001101110101110001001001111001;
		correct = 32'b01110010010011011000000000000000;
		#400 //4.070347e+30 * -451039000.0 = 4.070347e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100100000111101101000000100;
		b = 32'b10001010100100011000011101000111;
		correct = 32'b10010100100000111101101000001101;
		#400 //-1.3313612e-26 * -1.4013878e-32 = -1.3313626e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110101111010110100110110011;
		b = 32'b10010000000011111010000001110110;
		correct = 32'b00010110101111010110010100110110;
		#400 //3.0601302e-25 * -2.8325392e-29 = 3.059847e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011011111001111111001110001;
		b = 32'b11111001100111100000110111000100;
		correct = 32'b11111001100111100001010110101100;
		#400 //-2.0044243e+31 * -1.0258276e+35 = -1.0260281e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111110000100100000110001101;
		b = 32'b10010110001100110101010011100011;
		correct = 32'b11111111110000100100000110001101;
		#400 //nan * -1.448629e-25 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111001100110111110000110001;
		b = 32'b10101001100001011000101110111100;
		correct = 32'b11100111001100110111110000110001;
		#400 //-8.475945e+23 * -5.9306265e-14 = -8.475945e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010011100000100111110101001;
		b = 32'b00010111001000010110101100111110;
		correct = 32'b11001010011100000100111110101001;
		#400 //-3937258.2 * 5.2157264e-25 = -3937258.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101010010000101111000001101;
		b = 32'b10110000000010010101000011001011;
		correct = 32'b11011101010010000101111000001101;
		#400 //-9.023745e+17 * -4.9955123e-10 = -9.023745e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011001001110101011110110001110;
		b = 32'b00111011100110110101100011111001;
		correct = 32'b00111011100110110101100011111001;
		#400 //-9.654255e-24 * 0.004740831 = 0.004740831
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100011100001000001101001011;
		b = 32'b01111010110101100001011111100101;
		correct = 32'b01111010110101100001011111100101;
		#400 //-63049004.0 * 5.558181e+35 = 5.558181e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101101000111111000111101000;
		b = 32'b00010011100100001110110010000000;
		correct = 32'b01111101101000111111000111101000;
		#400 //2.7240027e+37 * 3.6583918e-27 = 2.7240027e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000110001001100111100111001;
		b = 32'b00000000100110111110110100010101;
		correct = 32'b00011000110001001100111100111001;
		#400 //5.0874054e-24 * 1.4319551e-38 = 5.0874054e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010001111110111110110011111;
		b = 32'b01110110011010110001011010110001;
		correct = 32'b01110110011010110001011010110000;
		#400 //-5.7874515e+25 * 1.192041e+33 = 1.1920409e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000011100100100011111110011;
		b = 32'b10001111101011101000100101100101;
		correct = 32'b01110000011100100100011111110011;
		#400 //2.9992941e+29 * -1.7210647e-29 = 2.9992941e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001011100100000111111111010;
		b = 32'b11011010010100001010100110110111;
		correct = 32'b11011010010100001010100110110111;
		#400 //-15.128901 * -1.468335e+16 = -1.468335e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001110111000001001010010111;
		b = 32'b00010010110101010101101110010101;
		correct = 32'b01100001110111000001001010010111;
		#400 //5.074529e+20 * 1.3464767e-27 = 5.074529e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010100110010001001110000101;
		b = 32'b00001001001101000000110000111110;
		correct = 32'b01000010100110010001001110000101;
		#400 //76.538124 * 2.1672468e-33 = 76.538124
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001010011101110001110010001;
		b = 32'b10010001011110111110011000100010;
		correct = 32'b10010001011110111110011011110001;
		#400 //-2.490335e-33 * -1.9871324e-28 = -1.9871573e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011000011010101101100001101;
		b = 32'b01111101101011011001101010100011;
		correct = 32'b01111101101011011001101010100011;
		#400 //-4.1540697e-37 * 2.884492e+37 = 2.884492e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111000011000101101110001011;
		b = 32'b11010110010100100100010110111011;
		correct = 32'b11100111000011000101101110001011;
		#400 //-6.6282e+23 * -57799233000000.0 = -6.6282e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110001000101101100111000001010;
		b = 32'b01101010001010100111010101110010;
		correct = 32'b01110001000101101101000010110100;
		#400 //7.467494e+29 * 5.1518e+25 = 7.468009e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101100001000100110110010101001;
		b = 32'b11110010111100010010100100010011;
		correct = 32'b11110010111100010010100100010011;
		#400 //2.3081903e-12 * -9.5533495e+30 = -9.5533495e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101010110110100101111100010;
		b = 32'b11011110011001001111100010101100;
		correct = 32'b11011110011001001111100010101100;
		#400 //-8.169428e-07 * -4.1247816e+18 = -4.1247816e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000100010010001101011001011;
		b = 32'b00000111111000100010110000011001;
		correct = 32'b00000111111000100010100111110101;
		#400 //-1.2591074e-38 * 3.403062e-34 = 3.402936e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111111110010010000000000000;
		b = 32'b10011101001000001110000101110110;
		correct = 32'b10111111111110010010000000000000;
		#400 //-1.9462891 * -2.1292384e-21 = -1.9462891
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000110111010011101101001111000;
		b = 32'b10000011101101011111000101110101;
		correct = 32'b10000110111011001011001000111110;
		#400 //-8.796587e-35 * -1.069366e-36 = -8.9035237e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101100000001101000110010010110;
		b = 32'b10000000001110111001100100111111;
		correct = 32'b00101100000001101000110010010110;
		#400 //1.9120586e-12 * -5.473269e-39 = 1.9120586e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001100100100010010000010000;
		b = 32'b10110111111010111010111110010100;
		correct = 32'b11000001100100100010010000011111;
		#400 //-18.267609 * -2.8095943e-05 = -18.267637
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011100110100101010010101111;
		b = 32'b00011100001000000100010010010101;
		correct = 32'b01101011100110100101010010101111;
		#400 //3.7314897e+26 * 5.30282e-22 = 3.7314897e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110001010000010110000000011;
		b = 32'b01101110011100101100111000110001;
		correct = 32'b01101110011100101100111000110001;
		#400 //-3.8237868e-11 * 1.8786161e+28 = 1.8786161e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000100001110010100000111111;
		b = 32'b10011110111101010001111111011101;
		correct = 32'b11000000100001110010100000111111;
		#400 //-4.223663 * -2.5953562e-20 = -4.223663
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010000110100001000100101111;
		b = 32'b00101001001000010100001001010001;
		correct = 32'b01001010000110100001000100101111;
		#400 //2524235.8 * 3.5806702e-14 = 2524235.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000000000100111110101010001;
		b = 32'b01000001011101010110011101011101;
		correct = 32'b11101000000000100111110101010001;
		#400 //-2.4648773e+24 * 15.337735 = -2.4648773e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011110010011110111101101011;
		b = 32'b10110001100101100010011010001001;
		correct = 32'b10110001100101100011001100101000;
		#400 //-1.4348361e-12 * -4.3699555e-09 = -4.3713904e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000010001001001010111001101;
		b = 32'b01011000110001011100110001001111;
		correct = 32'b01011000110001011100110001001111;
		#400 //-7.1517264e-10 * 1739850300000000.0 = 1739850300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001001101111001100011100010;
		b = 32'b00101101101001010100001011100101;
		correct = 32'b11111001001101111001100011100010;
		#400 //-5.9580697e+34 * 1.8788035e-11 = -5.9580697e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001111000010010100010010011;
		b = 32'b11001100100011010010101001100000;
		correct = 32'b01101001111000010010100010010011;
		#400 //3.402499e+25 * -74011390.0 = 3.402499e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100011110111111001010111101;
		b = 32'b00011100110000011011011100000000;
		correct = 32'b00011100110000011011011100000000;
		#400 //-1.9409383e-31 * 1.2818973e-21 = 1.2818973e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011100111100001110010111111;
		b = 32'b00011000111110001100111010000011;
		correct = 32'b01110011100111100001110010111111;
		#400 //2.5053892e+31 * 6.431502e-24 = 2.5053892e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110101001000011100101001000;
		b = 32'b00000101100001100000100100000111;
		correct = 32'b00101110101001000011100101001000;
		#400 //7.468032e-11 * 1.2604616e-35 = 7.468032e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100001110000011000100001010111;
		b = 32'b10111101000001001100111001010011;
		correct = 32'b10111101000001001100111001010011;
		#400 //-1.3114278e-18 * -0.03242333 = -0.03242333
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010100001111001101000000101;
		b = 32'b01000111100001100110111110001000;
		correct = 32'b01100010100001111001101000000101;
		#400 //1.2507044e+21 * 68831.06 = 1.2507044e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110111100010111010100101101;
		b = 32'b01111110111100010010101010111101;
		correct = 32'b01111110111100010010101010111101;
		#400 //7.1960008e-06 * 1.6028293e+38 = 1.6028293e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110100110000010001100110000100;
		b = 32'b00010000101011100010011000111001;
		correct = 32'b10110100110000010001100110000100;
		#400 //-3.5967616e-07 * 6.868979e-29 = -3.5967616e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110100111101010111010000011000;
		b = 32'b10000101001001111100001111101001;
		correct = 32'b10110100111101010111010000011000;
		#400 //-4.5719275e-07 * -7.888285e-36 = -4.5719275e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001010001011100011100000011;
		b = 32'b11010110100010111101001010000110;
		correct = 32'b11111001010001011100011100000011;
		#400 //-6.418243e+34 * -76868150000000.0 = -6.418243e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110100110000010001110010001;
		b = 32'b10100111111001101100111101010001;
		correct = 32'b10100111111001101100111101010001;
		#400 //2.457937e-25 * -6.4062597e-15 = -6.4062597e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110101000110101110111101111;
		b = 32'b01110000000110110101101010010011;
		correct = 32'b01110000000001101110111011010101;
		#400 //-2.5279808e+28 * 1.923187e+29 = 1.6703889e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110000100000100110111010100;
		b = 32'b10001111001100000001010100101111;
		correct = 32'b01010110000100000100110111010100;
		#400 //39665986000000.0 * -8.68155e-30 = 39665986000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001101001110101101111111000011;
		b = 32'b10111011011110110011001001111001;
		correct = 32'b10111011011110110011001001111001;
		#400 //-5.758502e-31 * -0.0038329645 = -0.0038329645
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110101100000000101000110011000;
		b = 32'b01101100001011100111000110000001;
		correct = 32'b11110101100000000101000110000010;
		#400 //-3.253266e+32 * 8.435564e+26 = -3.2532577e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010010000011100000110011100011;
		b = 32'b11100110110100101011000001110111;
		correct = 32'b11100110110100101011000001110111;
		#400 //-152525390000.0 * -4.9747608e+23 = -4.9747608e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111100001010100010110001101;
		b = 32'b11001001011110001110010001001001;
		correct = 32'b11001001011110001110010001001001;
		#400 //-3.6990323e-15 * -1019460.56 = -1019460.56
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111001010110011000110001111;
		b = 32'b01000100111001000000101111110010;
		correct = 32'b01000100111001000000101111110010;
		#400 //2.3757883e-15 * 1824.3733 = 1824.3733
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111100110111010110111111011;
		b = 32'b00110011101010101110110000010111;
		correct = 32'b10110111100110110000001100001111;
		#400 //-1.8558456e-05 * 7.9591864e-08 = -1.8478864e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011011011001100011111011111;
		b = 32'b11100111110101111111100110111101;
		correct = 32'b11100111110101111111100110111101;
		#400 //-6.9583607e-37 * -2.0398313e+24 = -2.0398313e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101111010010110010101101000;
		b = 32'b11000111000111111001000111010000;
		correct = 32'b11000111000111111001000111010000;
		#400 //4.0487773e-16 * -40849.812 = -40849.812
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100000110110011011010000010;
		b = 32'b01101001001010011110000100000100;
		correct = 32'b01101001001010011110000100000100;
		#400 //-7.83625e-27 * 1.2835692e+25 = 1.2835692e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000001100100100101011001111;
		b = 32'b11010110100111010100110111011100;
		correct = 32'b11010110100111010100110111011100;
		#400 //6.486233e-10 * -86478865000000.0 = -86478865000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010100110011110000111011110;
		b = 32'b10000000000000000001000100101001;
		correct = 32'b11110010100110011110000111011110;
		#400 //-6.0959057e+30 * -6.156e-42 = -6.0959057e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011100010001000010111000110;
		b = 32'b10100110000000111101011000000011;
		correct = 32'b11110011100010001000010111000110;
		#400 //-2.1632862e+31 * -4.5739795e-16 = -2.1632862e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100111111010101101101001000;
		b = 32'b10110001001000010010010100110101;
		correct = 32'b00111100111111010101101101000111;
		#400 //0.030927315 * -2.3449733e-09 = 0.030927313
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001000000101010101011101101;
		b = 32'b11001011110011010111011001011100;
		correct = 32'b11001011110011010111011001011100;
		#400 //1.0307862e-28 * -26930360.0 = -26930360.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001101001111000110011001000;
		b = 32'b11110010111110100100000101001100;
		correct = 32'b11110010111110100100000101001100;
		#400 //2.6434717e-28 * -9.9136245e+30 = -9.9136245e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111110010110100110110111000;
		b = 32'b01000101000111011111110110110110;
		correct = 32'b11011111110010110100110110111000;
		#400 //-2.9299135e+19 * 2527.857 = -2.9299135e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110001100010101000100110001;
		b = 32'b00100010111100110001001010000011;
		correct = 32'b11001110001100010101000100110001;
		#400 //-743722050.0 * 6.588488e-18 = -743722050.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101000110010100110101000001;
		b = 32'b10001011101100011000111111010010;
		correct = 32'b10011101000110010100110101000001;
		#400 //-2.028932e-21 * -6.8394317e-32 = -2.028932e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000100111001101110000001110;
		b = 32'b00011010111010101100010110100010;
		correct = 32'b00011010111010101100010110100010;
		#400 //-1.4405278e-38 * 9.7099425e-23 = 9.7099425e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001110011100000101100010100001;
		b = 32'b00011010101111101110001010000010;
		correct = 32'b01001110011100000101100010100001;
		#400 //1008085060.0 * 7.89481e-23 = 1008085060.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011100100110100010011111010;
		b = 32'b10110101101100000010100001001101;
		correct = 32'b10110101101100000010100001000100;
		#400 //1.0464123e-12 * -1.3124751e-06 = -1.3124741e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010010010010010110100001001;
		b = 32'b10010001110101101111111100101100;
		correct = 32'b01000010010010010010110100001001;
		#400 //50.29398 * -3.3920509e-28 = 50.29398
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100111010000100111101001000;
		b = 32'b10000101110001110010101011101110;
		correct = 32'b01110100111010000100111101001000;
		#400 //1.4724376e+32 * -1.872964e-35 = 1.4724376e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100001000011011110001010111;
		b = 32'b00001000000011001111001100101111;
		correct = 32'b11100100001000011011110001010111;
		#400 //-1.1933988e+22 * 4.241558e-34 = -1.1933988e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110010101110101011101000011;
		b = 32'b01100010001000100011001111110010;
		correct = 32'b01100010001000100011001111110010;
		#400 //-3.208829e-06 * 7.480289e+20 = 7.480289e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001111010010101000101010011;
		b = 32'b10000111111110001011110000101010;
		correct = 32'b11110001111010010101000101010011;
		#400 //-2.3106663e+30 * -3.7425486e-34 = -2.3106663e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001000110110010011000100000;
		b = 32'b11101001011110101110010100001010;
		correct = 32'b11101001011110101110010110100101;
		#400 //-1.7887453e+20 * -1.8957066e+25 = -1.8957245e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001000000111001011101010001;
		b = 32'b10110100001000101111010001011111;
		correct = 32'b10110100001000101111010001011111;
		#400 //4.458479e-19 * -1.5176327e-07 = -1.5176327e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001011010000001101000111011;
		b = 32'b10000011000111100111000000101010;
		correct = 32'b10110001011010000001101000111011;
		#400 //-3.3775354e-09 * -4.6560785e-37 = -3.3775354e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011111000110011100100101101;
		b = 32'b00111000111100000111111001100110;
		correct = 32'b01001011111000110011100100101101;
		#400 //29782618.0 * 0.00011467635 = 29782618.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110010111101001001101110110;
		b = 32'b11001011010010011110001110110101;
		correct = 32'b11001011010010011110001110110101;
		#400 //-5.0607928e-11 * -13231029.0 = -13231029.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101001111100000111111111001;
		b = 32'b10010010100111110001101100110010;
		correct = 32'b11010101001111100000111111111001;
		#400 //-13060988000000.0 * -1.0041015e-27 = -13060988000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011101110101010101011100101;
		b = 32'b10110010100101000011000111011010;
		correct = 32'b11111011101110101010101011100101;
		#400 //-1.9384667e+36 * -1.7252137e-08 = -1.9384667e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000110011011011111011010011;
		b = 32'b11110110010110111000101010011001;
		correct = 32'b11110110010110111010010001010001;
		#400 //-5.0940095e+29 * -1.1132071e+33 = -1.11371655e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111001100011101011001101111111;
		b = 32'b10000001111011100100100001011100;
		correct = 32'b00111001100011101011001101111111;
		#400 //0.00027218086 * -8.7531223e-38 = 0.00027218086
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111010100111100101011110011;
		b = 32'b11010010001101101110100000110100;
		correct = 32'b11010010001101101110100000110100;
		#400 //0.8273155 * -196394940000.0 = -196394940000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101101100011101000101011001;
		b = 32'b00111101011010000101101100011111;
		correct = 32'b11100101101100011101000101011001;
		#400 //-1.0496508e+23 * 0.056727525 = -1.0496508e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011110111100100111111100000001;
		b = 32'b10110111010000110000110001000111;
		correct = 32'b10110111010000110000110001000111;
		#400 //2.5675274e-20 * -1.1625764e-05 = -1.1625764e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010100001000000111000000110;
		b = 32'b00010110100001110000010011100101;
		correct = 32'b10111010100001000000111000000110;
		#400 //-0.001007498 * 2.1813515e-25 = -0.001007498
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110111010001111110010000110;
		b = 32'b00101110100000110111101011000010;
		correct = 32'b00111110111010001111110010000110;
		#400 //0.4550516 * 5.9789965e-11 = 0.4550516
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110011000011011010001110110;
		b = 32'b01000110101110011010110010111100;
		correct = 32'b01000111000101010100001101111100;
		#400 //14445.115 * 23766.367 = 38211.484
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100000101000010010010001110;
		b = 32'b01010011011001101101011011000010;
		correct = 32'b11111100000101000010010010001110;
		#400 //-3.0768054e+36 * 991445500000.0 = -3.0768054e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111100110011101000110010011;
		b = 32'b10000000101010101100001011110111;
		correct = 32'b11010111100110011101000110010011;
		#400 //-338250800000000.0 * -1.5681975e-38 = -338250800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111001101001001011011010111100;
		b = 32'b01111100011001110000100000011101;
		correct = 32'b01111100011001110000100000011101;
		#400 //0.00031416665 * 4.7983405e+36 = 4.7983405e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010101111011101011000000010001;
		b = 32'b11100011101011011100001111010110;
		correct = 32'b11100011101011011100001111010110;
		#400 //-9.640522e-26 * -6.4107964e+21 = -6.4107964e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001100111001001001000101111;
		b = 32'b10011011100101100101111011000110;
		correct = 32'b01100001100111001001001000101111;
		#400 //3.610282e+20 * -2.4876664e-22 = 3.610282e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011101111001111111001000010;
		b = 32'b11110100000010111000000111110011;
		correct = 32'b11110100000010111000000111110011;
		#400 //-4.770859e-27 * -4.421173e+31 = -4.421173e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100110100010000001110011111;
		b = 32'b10111010101010110011110010001000;
		correct = 32'b01110100110100010000001110011111;
		#400 //1.3247845e+32 * -0.0013064304 = 1.3247845e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000011100010000000001000010101;
		b = 32'b01100101111101011000001010000100;
		correct = 32'b01100101111101011000001010000100;
		#400 //7.99384e-37 * 1.4492342e+23 = 1.4492342e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101100100001001110010000000011;
		b = 32'b00000100011000011001100011100101;
		correct = 32'b10101100100001001110010000000011;
		#400 //-3.77698e-12 * 2.6518829e-36 = -3.77698e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011100101001010110010100100;
		b = 32'b10101001001011111111101100111100;
		correct = 32'b11101011100101001010110010100100;
		#400 //-3.594726e+26 * -3.9075717e-14 = -3.594726e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110111001010001111010110000100;
		b = 32'b11001101110110010100010100100001;
		correct = 32'b11110111001010001111010110000100;
		#400 //-3.4268966e+33 * -455648300.0 = -3.4268966e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111101001000010110100111010;
		b = 32'b01100101101001000011110110011011;
		correct = 32'b01100101101001000011110110011011;
		#400 //-4.556818e-15 * 9.6950565e+22 = 9.6950565e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101001010010011001010001100;
		b = 32'b10111110011110010011011101000000;
		correct = 32'b10111110011110010011011101000000;
		#400 //-7.955626e-36 * -0.24337482 = -0.24337482
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110010101001101100000110100;
		b = 32'b00010100100100111010110010111011;
		correct = 32'b00111110010101001101100000110100;
		#400 //0.207856 * 1.4911337e-26 = 0.207856
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110111100100011000110000111;
		b = 32'b00100011111011110110010100101101;
		correct = 32'b11010110111100100011000110000111;
		#400 //-133147270000000.0 * 2.5955282e-17 = -133147270000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110111110110010111001011010101;
		b = 32'b10011110011010010100001001010010;
		correct = 32'b01110111110110010111001011010101;
		#400 //8.8207616e+33 * -1.2348632e-20 = 8.8207616e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000001000100010011011110111;
		b = 32'b01101001011110111101010000101011;
		correct = 32'b01101001011110111101010000101011;
		#400 //-3.136385e-39 * 1.9027645e+25 = 1.9027645e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001100101101011010001011010;
		b = 32'b10010100000001001110001111110011;
		correct = 32'b00011001100101101010001110111110;
		#400 //1.558248e-23 * -6.709252e-27 = 1.5575771e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101011110101010000001111010;
		b = 32'b01000000111001110001000011110101;
		correct = 32'b01000000111001110001000011110101;
		#400 //1.17844184e-35 * 7.22082 = 7.22082
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001101001001100100110100110;
		b = 32'b11001110011001100100000100010000;
		correct = 32'b01010001101000101111110100100100;
		#400 //88469720000.0 * -965755900.0 = 87503960000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100000110100111000011011010;
		b = 32'b01001111100101000101110001100010;
		correct = 32'b01001111100101000101110001100010;
		#400 //-1.1897688e-31 * 4978164700.0 = 4978164700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110010011001000001010111001;
		b = 32'b10010101011111100010101001011111;
		correct = 32'b10101110010011001000001010111001;
		#400 //-4.6500335e-11 * -5.1328316e-26 = -4.6500335e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010000011001101111100010110;
		b = 32'b10000010001011000101001101111011;
		correct = 32'b11110010000011001101111100010110;
		#400 //-2.790246e+30 * -1.2660522e-37 = -2.790246e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011100100111110111111000110;
		b = 32'b00011111111000100110110010110110;
		correct = 32'b10101011100100111110111111000101;
		#400 //-1.0511529e-12 * 9.589457e-20 = -1.0511528e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001001010100100110000110111;
		b = 32'b00001100111111010000000110100001;
		correct = 32'b01101001001010100100110000110111;
		#400 //1.2867331e+25 * 3.8981802e-31 = 1.2867331e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010101100101100011111011110010;
		b = 32'b11000101101110110111110010100110;
		correct = 32'b11000101101110110111110010100110;
		#400 //6.068383e-26 * -5999.581 = -5999.581
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000000001101001111100001100101;
		b = 32'b00011100011010100000100000111011;
		correct = 32'b00011100011010100000100000111011;
		#400 //4.864553e-39 * 7.7434743e-22 = 7.7434743e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101001111111000010001110111;
		b = 32'b00000010111100101111001001011100;
		correct = 32'b10011101001111111000010001110111;
		#400 //-2.5347122e-21 * 3.5697812e-37 = -2.5347122e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101010100010001000100010101000;
		b = 32'b00010000100111111111000010111100;
		correct = 32'b00101010100010001000100010101000;
		#400 //2.4253277e-13 * 6.308535e-29 = 2.4253277e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100001010100000000001111100;
		b = 32'b10111010011110011001011111010001;
		correct = 32'b11110100001010100000000001111100;
		#400 //-5.387575e+31 * -0.00095212186 = -5.387575e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000101111110001010101111000;
		b = 32'b10001000010000001101010110101011;
		correct = 32'b01110000101111110001010101111000;
		#400 //4.7310073e+29 * -5.8029064e-34 = 4.7310073e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010101001111101011010001110;
		b = 32'b01000010100001110100010000000100;
		correct = 32'b01000010100001110100010000000100;
		#400 //-4.549261e-18 * 67.63284 = 67.63284
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000100011000001010110111000001;
		b = 32'b00000110010000010100101100001001;
		correct = 32'b00000110010011110101010111100101;
		#400 //2.6410857e-36 * 3.6354393e-35 = 3.8995478e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001001110111011011001010001;
		b = 32'b11000000011110111111101101110010;
		correct = 32'b11000001011110101011010100101110;
		#400 //-11.732011 * -3.937222 = -15.669233
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110110110011001100011000110;
		b = 32'b11110110011011101101100011011010;
		correct = 32'b11110110011011101101100011011010;
		#400 //-9.8951555e-11 * -1.21109856e+33 = -1.21109856e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101010101100011100100111011;
		b = 32'b10000110010101001101001011001100;
		correct = 32'b00110101010101100011100100111011;
		#400 //7.9804494e-07 * -4.0027637e-35 = 7.9804494e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110110001110100010111111101;
		b = 32'b00000111101101011000000111010101;
		correct = 32'b01000110110001110100010111111101;
		#400 //25506.994 * 2.7310162e-34 = 25506.994
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111001001100011000011111111100;
		b = 32'b11110100010111011111001001111100;
		correct = 32'b11110100010111011111001001111100;
		#400 //-0.00016930694 * -7.0337877e+31 = -7.0337877e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111100001101000111011101110;
		b = 32'b11011101011000001011000100010101;
		correct = 32'b11011111100011011001010001110111;
		#400 //-1.9391897e+19 * -1.0119216e+18 = -2.040382e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011101010110010001010001111;
		b = 32'b10110000100011101011100000101001;
		correct = 32'b10110000100011101011100000101001;
		#400 //1.8554493e-17 * -1.0384201e-09 = -1.0384201e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101110010000111001011011000;
		b = 32'b10001101111001010011010000101001;
		correct = 32'b11010101110010000111001011011000;
		#400 //-27549447000000.0 * -1.4125772e-30 = -27549447000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011110010101100010101011111;
		b = 32'b11111111010010010000101001000111;
		correct = 32'b11111111010010010000101001000111;
		#400 //-26577598.0 * -2.672282e+38 = -2.672282e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010001010000001111110010111;
		b = 32'b10100101111011111110100000101101;
		correct = 32'b11110010001010000001111110010111;
		#400 //-3.330027e+30 * -4.161722e-16 = -3.330027e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110100111110000111000110001101;
		b = 32'b00000001011111101010111100100001;
		correct = 32'b10110100111110000111000110001101;
		#400 //-4.627622e-07 * 4.677808e-38 = -4.627622e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110011010110110100111000010;
		b = 32'b10101011000001101001111010010101;
		correct = 32'b10110110011010110110100111000100;
		#400 //-3.5079288e-06 * -4.782644e-13 = -3.5079293e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000001101100010011101100011;
		b = 32'b00111000100111011000101110011000;
		correct = 32'b00111000100111011000101110011000;
		#400 //3.5923514e-29 * 7.512345e-05 = 7.512345e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000011111111101110100001111111;
		b = 32'b01110100001011010000011010111100;
		correct = 32'b01110100001011010000011010111100;
		#400 //1.4982157e-36 * 5.4834225e+31 = 5.4834225e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010001000000100011010011101;
		b = 32'b00001000101011001101110011010101;
		correct = 32'b10101010001000000100011010011101;
		#400 //-1.4235354e-13 * 1.0403791e-33 = -1.4235354e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100011101000001101101010110;
		b = 32'b00000110100000111000011100100000;
		correct = 32'b11101100011101000001101101010110;
		#400 //-1.18042796e+27 * 4.947527e-35 = -1.18042796e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100011001101101000011110001;
		b = 32'b00110000110000111010001001000110;
		correct = 32'b11101100011001101101000011110001;
		#400 //-1.11615855e+27 * 1.4234238e-09 = -1.11615855e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011100001110110110100110110;
		b = 32'b00111010100011100100101001001100;
		correct = 32'b11111011100001110110110100110110;
		#400 //-1.4063503e+36 * 0.0010855882 = -1.4063503e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011100111100110110000011001;
		b = 32'b00011110111101001100101000010100;
		correct = 32'b01111011100111100110110000011001;
		#400 //1.6451508e+36 * 2.5918082e-20 = 1.6451508e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001101011110110011110000010;
		b = 32'b10111100110011101001111001000000;
		correct = 32'b11011001101011110110011110000010;
		#400 //-6171491000000000.0 * -0.025221944 = -6171491000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100000011101010100111011010;
		b = 32'b01000101010000100000001001000000;
		correct = 32'b11101100000011101010100111011010;
		#400 //-6.898783e+26 * 3104.1406 = -6.898783e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001001110101011011001101010;
		b = 32'b01100001101101101010101101001111;
		correct = 32'b01100001101101101010101101001111;
		#400 //50120270000.0 * 4.2120644e+20 = 4.2120644e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010100001011100111100000101;
		b = 32'b11010100111000111110000000001100;
		correct = 32'b01101010100001011100111100000101;
		#400 //8.088238e+25 * -7829731700000.0 = 8.088238e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011111101111011011110100111;
		b = 32'b01110100100110001000110100010111;
		correct = 32'b01110100100110001000110100010111;
		#400 //-1.455952e-36 * 9.669077e+31 = 9.669077e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100010010000010001111111110;
		b = 32'b01000110101101110111010011111000;
		correct = 32'b11110100010010000010001111111110;
		#400 //-6.3427086e+31 * 23482.484 = -6.3427086e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011000011000011001001000101;
		b = 32'b00100100100010101001101111000011;
		correct = 32'b00100100100010101001101111000011;
		#400 //1.769527e-27 * 6.011183e-17 = 6.011183e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100010000110100010011111010;
		b = 32'b11110111010011110011001110000111;
		correct = 32'b11110111010011110011001110000111;
		#400 //-6.460924e-22 * -4.2025412e+33 = -4.2025412e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010000100101100010011011011;
		b = 32'b10100100110100101110100101011101;
		correct = 32'b10101010000100101101111100111000;
		#400 //-1.3035703e-13 * -9.1468315e-17 = -1.304485e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100010011001011110000100000101;
		b = 32'b00100000101100100100111011000001;
		correct = 32'b11100010011001011110000100000101;
		#400 //-1.0601297e+21 * 3.0206488e-19 = -1.0601297e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111000011001110100001100111;
		b = 32'b01010001001011001010000011100010;
		correct = 32'b01010111000011001111001100110001;
		#400 //154929790000000.0 * 46339596000.0 = 154976130000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001111000111010000100011100;
		b = 32'b11101000110101111000001110001011;
		correct = 32'b11101000110101110111111111111100;
		#400 //5.248775e+20 * -8.1418827e+24 = -8.1413575e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001110111111101010111110111;
		b = 32'b10000011101111010100100001000001;
		correct = 32'b11010001110111111101010111110111;
		#400 //-120170930000.0 * -1.112501e-36 = -120170930000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110010111101011100111101100;
		b = 32'b00010100100110001000110111011110;
		correct = 32'b10110110010111101011100111101100;
		#400 //-3.3188799e-06 * 1.5404035e-26 = -3.3188799e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111001011011001000101101000001;
		b = 32'b10110010001011101000011011011011;
		correct = 32'b00111001011011001000100010000111;
		#400 //0.0002255859 * -1.0158796e-08 = 0.00022557574
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001101001001010001111100100110;
		b = 32'b11110110110111011101110000100000;
		correct = 32'b11110110110111011101110000100000;
		#400 //-5.0882044e-31 * -2.2499263e+33 = -2.2499263e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111010101011101010100010000;
		b = 32'b11100100011000001110101110011000;
		correct = 32'b11100100011000001110101110011000;
		#400 //2.967519e-15 * -1.6596188e+22 = -1.6596188e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010000011001001110111000011;
		b = 32'b11111001010010001111010010110100;
		correct = 32'b11111001010010001111010010110100;
		#400 //-1.2489232e-13 * -6.521391e+34 = -6.521391e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101000001011010111100101000;
		b = 32'b10001000001111111101000101010100;
		correct = 32'b11000101000001011010111100101000;
		#400 //-2138.9473 * -5.7723036e-34 = -2138.9473
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011011010111101110010110010;
		b = 32'b10101011111101010011110001101110;
		correct = 32'b01011011011010111101110010110010;
		#400 //6.6389277e+16 * -1.742507e-12 = 6.6389277e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111100011011010100110101000;
		b = 32'b10111100110101011100010000110100;
		correct = 32'b00111111100010100101001010010111;
		#400 //1.10674 * -0.026094534 = 1.0806454
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110010000000011110100111111;
		b = 32'b11001100100000000011110000011110;
		correct = 32'b11001100100000000011110000011110;
		#400 //-4.3710143e-11 * -67231980.0 = -67231980.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101011011101110101000001011;
		b = 32'b10001010001111110100001111001111;
		correct = 32'b00011101011011101110101000001011;
		#400 //3.1620035e-21 * -9.209069e-33 = 3.1620035e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011001001111110011101000100001;
		b = 32'b11001100101011000000010101100101;
		correct = 32'b11001100101011000000010101100101;
		#400 //-9.8862076e-24 * -90188584.0 = -90188584.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100100100100111101010011110;
		b = 32'b10001010100100011101100101011011;
		correct = 32'b01101100100100100111101010011110;
		#400 //1.4166577e+27 * -1.4044752e-32 = 1.4166577e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101000001001010100110101011;
		b = 32'b01001001100010100110111000111101;
		correct = 32'b11100101000001001010100110101011;
		#400 //-3.9155137e+22 * 1134023.6 = -3.9155137e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111100100111111110100011101;
		b = 32'b11101001111011100100011100000111;
		correct = 32'b11101001111011100100011100000111;
		#400 //6.267566e-20 * -3.600747e+25 = -3.600747e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100001001011110111010011011;
		b = 32'b00000101011011100110010110110001;
		correct = 32'b00001100001001011111001001010101;
		#400 //1.278294e-31 * 1.1209384e-35 = 1.2784062e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111001000011111111110111111;
		b = 32'b01001101011101110011000100100101;
		correct = 32'b01001101011101110011000100100101;
		#400 //9.655893e-06 * 259199570.0 = 259199570.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101101001010011101100101001;
		b = 32'b01010000100001111101000011001110;
		correct = 32'b01010000100001111101000011001110;
		#400 //-1.87846e-11 * 18228867000.0 = 18228867000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010011101000010001001000010;
		b = 32'b10010100110010011100000010011111;
		correct = 32'b10010100110100010110000110110001;
		#400 //-7.703505e-28 * -2.0371789e-26 = -2.114214e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110110010010011000010100001;
		b = 32'b01010000100111111100011111101010;
		correct = 32'b01010000100111111100011111101010;
		#400 //7.567925e-35 * 21445431000.0 = 21445431000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011110001011010100110000111;
		b = 32'b10011011110100000100110011111010;
		correct = 32'b01000011110001011010100110000111;
		#400 //395.32443 * -3.4460458e-22 = 395.32443
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011000001111010010111100010;
		b = 32'b01110000010100101110111001010011;
		correct = 32'b01111011000001111010010111100101;
		#400 //7.043246e+35 * 2.6111987e+29 = 7.043248e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100110000001000011011011101;
		b = 32'b01001101110010110110110010100111;
		correct = 32'b11110100110000001000011011011101;
		#400 //-1.2202836e+32 * 426611940.0 = -1.2202836e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100111011100101101001111111;
		b = 32'b01111001011111001000000010101111;
		correct = 32'b01111001011111001000000010101111;
		#400 //-1.5772912e-21 * 8.19418e+34 = 8.19418e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111010011010011011010110100;
		b = 32'b00101000010111110010000110001001;
		correct = 32'b01001111010011010011011010110100;
		#400 //3442914300.0 * 1.23862585e-14 = 3442914300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001010000110000101100111010;
		b = 32'b00100110101101010100011100000000;
		correct = 32'b00100110101101010100011100000000;
		#400 //-3.5823898e-38 * 1.2578643e-15 = 1.2578643e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000101011111000000010011111;
		b = 32'b10101100101100101000100010010000;
		correct = 32'b10101100101100101000100010010000;
		#400 //1.0562668e-33 * -5.0742258e-12 = -5.0742258e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111110011001011000010101100;
		b = 32'b11100001011101000100101100011100;
		correct = 32'b11100001011101000100101100011100;
		#400 //6868261000.0 * -2.8165111e+20 = -2.8165111e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101100110010100010000001110011;
		b = 32'b11111000001001110100001010111101;
		correct = 32'b11111000001001110100001010111101;
		#400 //5.744788e-12 * -1.35698e+34 = -1.35698e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111101001110010010010111111;
		b = 32'b11000011101010110110100001101011;
		correct = 32'b01001111101001110010010010111110;
		#400 //5608406500.0 * -342.81577 = 5608406000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000110001001110011000011100;
		b = 32'b01101101101010101011011001101000;
		correct = 32'b01101101101010101011011001101000;
		#400 //26427318000.0 * 6.604121e+27 = 6.604121e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101000110001100111001101011;
		b = 32'b11111101000000001001001100110000;
		correct = 32'b11111101000000001001001100110000;
		#400 //-1.3253836e-16 * -1.0681589e+37 = -1.0681589e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111011011110100011010000010;
		b = 32'b10011100101110010100101101101101;
		correct = 32'b11111111011011110100011010000010;
		#400 //-3.1805159e+38 * -1.226177e-21 = -3.1805159e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010011001111110100001101111;
		b = 32'b00001111011110100001101110010000;
		correct = 32'b00001111011110100101010110001010;
		#400 //1.1165961e-32 * 1.233126e-29 = 1.2342426e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001101010001100000110000111;
		b = 32'b01001000001110010011100100011100;
		correct = 32'b01001000001110010011100100011100;
		#400 //1.7448958e-23 * 189668.44 = 189668.44
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000000010101000110001011011;
		b = 32'b11010101001010000101001100101011;
		correct = 32'b11011000000011010010110110101000;
		#400 //-609341700000000.0 * -11567197000000.0 = -620908900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010001010100101001101010100;
		b = 32'b11000011110110101100010010001010;
		correct = 32'b11000011110110101100010010001010;
		#400 //3.5222488e-23 * -437.53546 = -437.53546
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110100101111100111010100001;
		b = 32'b01100010011110001001101101101000;
		correct = 32'b11101110100101111100111010100001;
		#400 //-2.3491018e+28 * 1.1464977e+21 = -2.3491018e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100000010000011110001100111;
		b = 32'b11101011111001000010110010101101;
		correct = 32'b11111100000010000011110001100111;
		#400 //-2.82951e+36 * -5.5169212e+26 = -2.82951e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110001011101101001011111011;
		b = 32'b01011011001100010010111010010101;
		correct = 32'b11100110001011101101001011111000;
		#400 //-2.0639592e+23 * 4.987229e+16 = -2.0639586e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100001000111101011110000100;
		b = 32'b11101011110000111111010010011000;
		correct = 32'b01111100001000111101011110000100;
		#400 //3.4028623e+36 * -4.737912e+26 = 3.4028623e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111110010100111000100001100;
		b = 32'b11011100011110100001001010101000;
		correct = 32'b11011100011110100001001010101000;
		#400 //-1.9962282e-29 * -2.8155703e+17 = -2.8155703e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000000001001011011100010110100;
		b = 32'b01011000101000100000110101000011;
		correct = 32'b01011000101000100000110101000011;
		#400 //3.464172e-39 * 1425422700000000.0 = 1425422700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000101110011011010000100000;
		b = 32'b11011010001100011010110011001011;
		correct = 32'b11011010001100011010110011001011;
		#400 //1.117663e-33 * -1.2502765e+16 = -1.2502765e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001000010100100000111101100;
		b = 32'b00110000100001000111111101110110;
		correct = 32'b11011001000010100100000111101100;
		#400 //-2432251800000000.0 * 9.640491e-10 = -2432251800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011111100010110110000010000;
		b = 32'b11001000110111110000001101000001;
		correct = 32'b11001011111101001110100000011101;
		#400 //-31643680.0 * -456730.03 = -32100410.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111000010010110000100100110;
		b = 32'b01010010011110010111101011110100;
		correct = 32'b01010010011101110101010101101111;
		#400 //-2304845300.0 * 267877420000.0 = 265572560000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111010111110010011110110001;
		b = 32'b10000100000000001111111111110110;
		correct = 32'b00100111010111110010011110110001;
		#400 //3.0968984e-15 * -1.516386e-36 = 3.0968984e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010001000011001101001010001;
		b = 32'b10111101110101001100001100010011;
		correct = 32'b11101010001000011001101001010001;
		#400 //-4.884145e+25 * -0.1038877 = -4.884145e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110111010000010001000001101;
		b = 32'b10100111011000111010101111010000;
		correct = 32'b00101110111010000010000001000110;
		#400 //1.0556187e-10 * -3.1595718e-15 = 1.05558715e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000001101101001111010011000100;
		b = 32'b00010101000010110110110111010000;
		correct = 32'b00010101000010110110110111010000;
		#400 //6.647278e-38 * 2.8157453e-26 = 2.8157453e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010011000001100011101101110;
		b = 32'b11001000110110101001111000000011;
		correct = 32'b01100010011000001100011101101110;
		#400 //1.0366103e+21 * -447728.1 = 1.0366103e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011001111000010101011101100;
		b = 32'b10111101101010110100110100100110;
		correct = 32'b01100011001111000010101011101100;
		#400 //3.4710807e+21 * -0.08364324 = 3.4710807e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001001001100100011100100001;
		b = 32'b11111000100100100101001100011011;
		correct = 32'b11111000100100100101001100011011;
		#400 //8.596363e-24 * -2.374253e+34 = -2.374253e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000100011101001110100011010;
		b = 32'b00110000100010000111001011011111;
		correct = 32'b01001000100011101001110100011010;
		#400 //292072.8 * 9.927951e-10 = 292072.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010101110100100110011011001001;
		b = 32'b11101010101000000111101111001111;
		correct = 32'b11101010101000000111101111001111;
		#400 //-8.498049e-26 * -9.70064e+25 = -9.70064e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100111101111001110101101011;
		b = 32'b10111010111101000011001110110101;
		correct = 32'b01100100111101111001110101101011;
		#400 //3.6541512e+22 * -0.0018631133 = 3.6541512e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100000101011110010011000100011;
		b = 32'b10010001010101100101010111000010;
		correct = 32'b11100000101011110010011000100011;
		#400 //-1.0096651e+20 * -1.690805e-28 = -1.0096651e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100101111111100111101001100;
		b = 32'b00101011000000001110011010001111;
		correct = 32'b11111100101111111100111101001100;
		#400 //-7.9674654e+36 * 4.57947e-13 = -7.9674654e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101101001100000100100110101100;
		b = 32'b10010000011001001010011100001001;
		correct = 32'b00101101001100000100100110101100;
		#400 //1.00208e-11 * -4.509375e-29 = 1.00208e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111000110101110011101011000;
		b = 32'b10011010110001001100010001010011;
		correct = 32'b11101111000110101110011101011000;
		#400 //-4.794037e+28 * -8.138088e-23 = -4.794037e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101111011111100011010100111;
		b = 32'b11100110001110111100000101110010;
		correct = 32'b11100110001110111100000101110010;
		#400 //1.7864703e-06 * -2.2166274e+23 = -2.2166274e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100101000101001110011010000;
		b = 32'b01000010010001100111010111101001;
		correct = 32'b01000100101010001101000001111111;
		#400 //1300.9004 * 49.615147 = 1350.5155
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100010100111111110110001000;
		b = 32'b01111000110111000000010000100110;
		correct = 32'b01111100010101011011010110010000;
		#400 //4.4028674e+36 * 3.569967e+34 = 4.438567e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111000010000111000000011100;
		b = 32'b11110001110011001100111101001001;
		correct = 32'b11110001110011001100111101001001;
		#400 //34928.11 * -2.0283371e+30 = -2.0283371e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001001011011101000010010011;
		b = 32'b01101000010000010111110010001000;
		correct = 32'b01101000010000010111110010001000;
		#400 //3.8594626e-14 * 3.6548557e+24 = 3.6548557e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100110100100010111100001111;
		b = 32'b10001101011101011011110011001001;
		correct = 32'b01101100110100100010111100001111;
		#400 //2.0327732e+27 * -7.5723696e-31 = 2.0327732e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010010111111110010000110100;
		b = 32'b00110111111001010101001011100001;
		correct = 32'b00110111111001010101001011100001;
		#400 //-1.077998e-32 * 2.733752e-05 = 2.733752e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101000011101011101000001000;
		b = 32'b10001100010000111001101100001000;
		correct = 32'b11001101000011101011101000001000;
		#400 //-149659780.0 * -1.5068907e-31 = -149659780.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111000011111110110101111001;
		b = 32'b01111001111110100011110110000100;
		correct = 32'b01111001111110100011110110000100;
		#400 //6.79679e+23 * 1.6241524e+35 = 1.6241524e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011000111000010101010111111;
		b = 32'b11100000010011101001010100101001;
		correct = 32'b11100011000111110110010100010100;
		#400 //-2.8807723e+21 * -5.9543397e+19 = -2.9403158e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000001110100100100000101111;
		b = 32'b01011101100010010001000110011000;
		correct = 32'b01100000001111101001000010111100;
		#400 //5.369212e+19 * 1.2346053e+18 = 5.492673e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110100000000011001100000101;
		b = 32'b11011010000110110110101111000110;
		correct = 32'b11011010000110110110101111000110;
		#400 //-3.1603566e-30 * -1.093678e+16 = -1.093678e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011000001010011011001011011;
		b = 32'b01111101011000010110000111100101;
		correct = 32'b01111101011000010110000111100101;
		#400 //-0.0020326588 * 1.8724037e+37 = 1.8724037e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100011000001000110111100000110;
		b = 32'b01101010101110001000010101011111;
		correct = 32'b01101010101110001000010101011111;
		#400 //-7.1792445e-18 * 1.1153609e+26 = 1.1153609e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101100000000101001111110010;
		b = 32'b00001101100110001011011001001010;
		correct = 32'b00011101100000000101001111110010;
		#400 //3.3968115e-21 * 9.411608e-31 = 3.3968115e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000000000100110101011000100;
		b = 32'b11101001111000010010100010010101;
		correct = 32'b11101001111000010010100010000101;
		#400 //3.7590156e+19 * -3.4024994e+25 = -3.4024957e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111110111101010011111010010;
		b = 32'b10000111011111011101000010011001;
		correct = 32'b00001111110111101010011101010011;
		#400 //2.1955532e-29 * -1.9094906e-34 = 2.1955341e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100100011110110000001010101;
		b = 32'b10100110010110000000110001110000;
		correct = 32'b11011100100011110110000001010101;
		#400 //-3.2285472e+17 * -7.495691e-16 = -3.2285472e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110111011111111110001011110;
		b = 32'b10011111001111111000100001000010;
		correct = 32'b11010110111011111111110001011110;
		#400 //-131933590000000.0 * -4.0558533e-20 = -131933590000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111010100111111001100000100;
		b = 32'b10101010000001011100000001100111;
		correct = 32'b10110111010100111111001100000100;
		#400 //-1.26331615e-05 * -1.1879526e-13 = -1.26331615e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100111110101000100111100001;
		b = 32'b11100110111001101110000100110001;
		correct = 32'b11100110111001101110000100110001;
		#400 //-131354376.0 * -5.4514917e+23 = -5.4514917e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101010011111010011110000000;
		b = 32'b01100101100100010000111010101100;
		correct = 32'b01100101100100010000111010101100;
		#400 //-0.05069685 * 8.562672e+22 = 8.562672e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101011101101101100111001100;
		b = 32'b11010100110011110111000010000101;
		correct = 32'b11010100110011110111000010000101;
		#400 //1.16068674e-35 * -7127568000000.0 = -7127568000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111011010001110111010111001;
		b = 32'b01111000011101101011101001100000;
		correct = 32'b01111000011101101011101001100000;
		#400 //-1.6784556e+19 * 2.0016956e+34 = 2.0016956e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011111110011101000110001101;
		b = 32'b10011101010111000101001101000100;
		correct = 32'b10011101010111000101001101000100;
		#400 //-1.4683015e-36 * -2.9159805e-21 = -2.9159805e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000000111110100101100111110;
		b = 32'b00011111111100000110010110101000;
		correct = 32'b00011111111100000110010110101000;
		#400 //3.1415185e-29 * 1.0181213e-19 = 1.0181213e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110111101011110100100000100;
		b = 32'b11110101100000011100010101111101;
		correct = 32'b11111110111101011110100100100100;
		#400 //-1.6343537e+38 * -3.290097e+32 = -1.634357e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011110000010010000111101111;
		b = 32'b11100101111000011000011011010010;
		correct = 32'b11100101111000011000011011011110;
		#400 //-1.0872396e+17 * -1.3312743e+23 = -1.3312754e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110110000110010100110110011;
		b = 32'b11011010001111010000111110011001;
		correct = 32'b11011010001111010000111110011001;
		#400 //-5.8163073e-06 * -1.330398e+16 = -1.330398e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001101001100111101111000100;
		b = 32'b01101001111001011111001010111110;
		correct = 32'b01101001111001011111001010111110;
		#400 //1.1281358e-18 * 3.4748791e+25 = 3.4748791e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110100101100000110011101000;
		b = 32'b01100011011010110100010101100100;
		correct = 32'b11111110100101100000110011101000;
		#400 //-9.972561e+37 * 4.339985e+21 = -9.972561e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001010100110010101111110101;
		b = 32'b01010100100110000111101010001110;
		correct = 32'b11110001010100110010101111110101;
		#400 //-1.04567165e+30 * 5239129000000.0 = -1.04567165e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100011110110101101000111011;
		b = 32'b01000111101000101000110000100110;
		correct = 32'b01000111101001001000001011011010;
		#400 //1005.40985 * 83224.3 = 84229.7
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101011101111011101101001000;
		b = 32'b11100010011101110001000110110011;
		correct = 32'b11100010011101110001000110110011;
		#400 //17023984000000.0 * -1.1394053e+21 = -1.1394053e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011110100111110000101100011100;
		b = 32'b11001100100100010111010111001011;
		correct = 32'b11001100100100010111010111001011;
		#400 //1.6839375e-20 * -76263000.0 = -76263000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101000101000001001100100011;
		b = 32'b11101110100000001010110011011000;
		correct = 32'b01111101000101000001001100100011;
		#400 //1.2301569e+37 * -1.9911518e+28 = 1.2301569e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100110000001110000010011100;
		b = 32'b10011111000111111000001101011100;
		correct = 32'b00111100110000001110000010011100;
		#400 //0.023544602 * -3.3778218e-20 = 0.023544602
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100101010000101001111010010;
		b = 32'b00100101000001101001110100000010;
		correct = 32'b00110100101010000101001111010010;
		#400 //3.1353426e-07 * 1.1675844e-16 = 3.1353426e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011101110000101101001010110;
		b = 32'b10100001111011000001001111010111;
		correct = 32'b11011011101110000101101001010110;
		#400 //-1.0378144e+17 * -1.5997234e-18 = -1.0378144e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000011000011111011010101000100;
		b = 32'b00100010011011001111000000000001;
		correct = 32'b00100010011011001111000000000001;
		#400 //4.2232006e-37 * 3.2111021e-18 = 3.2111021e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110110101100111000010101000000;
		b = 32'b10001000110100101001110000111001;
		correct = 32'b01110110101100111000010101000000;
		#400 //1.8205542e+33 * -1.2675643e-33 = 1.8205542e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001001111110100010010101110;
		b = 32'b00010111011001001001000101110001;
		correct = 32'b00010111011001001001000101110001;
		#400 //2.3023082e-33 * 7.3854346e-25 = 7.3854346e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010010110001001010101010000110;
		b = 32'b01011000100010000100110111101011;
		correct = 32'b01011000100010000100000110100000;
		#400 //-422337250000.0 * 1198945900000000.0 = 1198523500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010111010110010101000101111;
		b = 32'b00010010010000000101001100010001;
		correct = 32'b00011010111010110010101010001111;
		#400 //9.7261873e-23 * 6.0686905e-28 = 9.726248e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111000110011001001101101011111;
		b = 32'b11010110011101101010100101001000;
		correct = 32'b11010110011101101010100101001000;
		#400 //9.756418e-05 * -67801730000000.0 = -67801730000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111101110100111101000101111;
		b = 32'b01100010001101001100010101110011;
		correct = 32'b01100010001110101001100101000100;
		#400 //2.6874208e+19 * 8.336604e+20 = 8.605346e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000010011100011010100010000;
		b = 32'b01010101111111110100001100111011;
		correct = 32'b01010101111111110100001100111011;
		#400 //211156.25 * 35083027000000.0 = 35083027000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001111011100100110111111100;
		b = 32'b10110001010010000111101110110011;
		correct = 32'b01001001111011100100110111111100;
		#400 //1952191.5 * -2.9174145e-09 = 1952191.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100010100110000010101101000;
		b = 32'b11010100011101000110100101101111;
		correct = 32'b11010100111000111011011101101100;
		#400 //-3625315200000.0 * -4198963600000.0 = -7824279000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001111101100011110111101111;
		b = 32'b00110011000110010100101001111110;
		correct = 32'b11001001111101100011110111101111;
		#400 //-2017213.9 * 3.569084e-08 = -2017213.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111000000000000100110000011;
		b = 32'b10101101011111011011011001010011;
		correct = 32'b11010111000000000000100110000011;
		#400 //-140778340000000.0 * -1.4421869e-11 = -140778340000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011011010000001100000111011;
		b = 32'b00100010100000100100001010000110;
		correct = 32'b11111011011010000001100000111011;
		#400 //-1.2051043e+36 * 3.5307005e-18 = -1.2051043e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001001100110011101111000100;
		b = 32'b11101110111111000001111001000100;
		correct = 32'b11101110111111000001111001000100;
		#400 //9.266153e-24 * -3.9013406e+28 = -3.9013406e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101000010011001010000110001;
		b = 32'b11101011011110110000110000110101;
		correct = 32'b11101011011110110000110000110101;
		#400 //-6.1960016e+17 * -3.0349803e+26 = -3.0349803e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100100001101001001010000101;
		b = 32'b10100100110000001110000001010000;
		correct = 32'b10111100100001101001001010000101;
		#400 //-0.016427288 * -8.364673e-17 = -0.016427288
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011111110100010010010111000;
		b = 32'b11011100111100011011001111001101;
		correct = 32'b11011100111100011011001111001101;
		#400 //-1.470211e-36 * -5.442653e+17 = -5.442653e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111111110011101000000000111;
		b = 32'b11010110101010011011000000111110;
		correct = 32'b11101111111110011101000000000111;
		#400 //-1.5462651e+29 * -93287210000000.0 = -1.5462651e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110001110101100001011000011;
		b = 32'b00001011100101001101010111010000;
		correct = 32'b01011110001110101100001011000011;
		#400 //3.3643833e+18 * 5.7329236e-32 = 3.3643833e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100111011011010100110000111;
		b = 32'b11010101011110110000101001100100;
		correct = 32'b01101100111011011010100110000111;
		#400 //2.2985279e+27 * -17251378000000.0 = 2.2985279e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011001001100111011000110110;
		b = 32'b00101111111011000100001110110000;
		correct = 32'b11111011001001100111011000110110;
		#400 //-8.643189e+35 * 4.2976245e-10 = -8.643189e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110101001000100011100110010;
		b = 32'b11010001101011110001011101101100;
		correct = 32'b11010001101011110001011101101100;
		#400 //2.654056e-25 * -94001530000.0 = -94001530000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101011011110001101011101110;
		b = 32'b01001100111100011010100100101101;
		correct = 32'b01001100111100011010100100101101;
		#400 //2.073907e-16 * 126699880.0 = 126699880.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110110100111101001101110000;
		b = 32'b11101101011010001010100110001101;
		correct = 32'b11101101011010001010100110001101;
		#400 //7.968006e-35 * -4.5003435e+27 = -4.5003435e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001101110100111111011001001;
		b = 32'b11111000000110100001000111011010;
		correct = 32'b11111000000110100001000111011010;
		#400 //1.263741e-18 * -1.2499622e+34 = -1.2499622e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011000011011010111110011011;
		b = 32'b11001100011010010000101100111000;
		correct = 32'b01110011000011011010111110011011;
		#400 //1.1225518e+31 * -61091040.0 = 1.1225518e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010111001101111111001100111;
		b = 32'b01111011111101011010000111111100;
		correct = 32'b01111011111101011010000111111100;
		#400 //6.2610984e-18 * 2.5507963e+36 = 2.5507963e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110110011110111000010001010;
		b = 32'b00010111010010000101011010001100;
		correct = 32'b11111110110011110111000010001010;
		#400 //-1.3786727e+38 * 6.4732723e-25 = -1.3786727e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111101100101001110010110111;
		b = 32'b00111001011000001001001110000010;
		correct = 32'b00111001011101101110011100011001;
		#400 //2.129223e-05 * 0.00021417256 = 0.00023546479
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101101000100000111101110010;
		b = 32'b01101011001111010100101110001000;
		correct = 32'b01101101101001111111100111001110;
		#400 //6.2694055e+27 * 2.2884367e+26 = 6.498249e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000011101111011110110110000;
		b = 32'b01001100101010101010000000110001;
		correct = 32'b01001100101010101010000000110001;
		#400 //4.885829e-29 * 89457030.0 = 89457030.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100100100110011110111001000;
		b = 32'b10101001110110101101100010001011;
		correct = 32'b10101001110110101101100010001011;
		#400 //-9.743614e-22 * -9.718709e-14 = -9.718709e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000011111011110000011101111;
		b = 32'b00110010101001010110000001010010;
		correct = 32'b01001000011111011110000011101111;
		#400 //259971.73 * 1.925233e-08 = 259971.73
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000101011010111101001001000;
		b = 32'b11100110010111000011010110110011;
		correct = 32'b11100110010111000011010110110011;
		#400 //6.842487e-29 * -2.599778e+23 = -2.599778e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100000101010111100101011011;
		b = 32'b00100101011101110111000010101001;
		correct = 32'b01011100000101010111100101011011;
		#400 //1.6829281e+17 * 2.1462006e-16 = 1.6829281e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111000000011110000110000010;
		b = 32'b10000001111101010000011000011010;
		correct = 32'b00111111000000011110000110000010;
		#400 //0.5073472 * -9.000754e-38 = 0.5073472
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101110000001010100000000010;
		b = 32'b11101010101011010100100001011101;
		correct = 32'b11101010101011010100100001011101;
		#400 //-1.811731e-35 * -1.0474295e+26 = -1.0474295e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110010010111010011010000000;
		b = 32'b00100001111111010010011111000110;
		correct = 32'b01010110010010111010011010000000;
		#400 //55978993000000.0 * 1.7154475e-18 = 55978993000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000000101101100011001111111;
		b = 32'b01010101011001000110000100001010;
		correct = 32'b01010101011001000110000100001010;
		#400 //-2.97352e-29 * 15694089000000.0 = 15694089000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011110100011000101001111101;
		b = 32'b11000001010101000111111011010101;
		correct = 32'b11000001010101000111111011010101;
		#400 //-9.757512e-08 * -13.280965 = -13.280965
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111000111101110001110011010;
		b = 32'b01010111000010101111011110010001;
		correct = 32'b01100111000111101110001110011010;
		#400 //7.503324e+23 * 152795900000000.0 = 7.503324e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001101101111001100000011000;
		b = 32'b00100100011101011110011110101001;
		correct = 32'b00101001101101111011011011010101;
		#400 //8.1532166e-14 * 5.332213e-17 = 8.158549e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100011101000101101101111101011;
		b = 32'b11110011110100000011001111111000;
		correct = 32'b11110011110100000011001111111000;
		#400 //-1.7657214e-17 * -3.2991083e+31 = -3.2991083e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111110101101100110110001111;
		b = 32'b11101110000111110110010110101011;
		correct = 32'b01111111110101101100110110001111;
		#400 //nan * -1.2332756e+28 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011110011111110001100010101;
		b = 32'b00011010101011111011011011100101;
		correct = 32'b00111011110011111110001100010101;
		#400 //0.006344209 * 7.2673786e-23 = 0.006344209
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011110111001010100101010010;
		b = 32'b01001111000010011000101101011000;
		correct = 32'b01001111000010011000101101011000;
		#400 //2.3924158e-17 * 2307610600.0 = 2307610600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000001000011100101100110011;
		b = 32'b11101101010100111101110101101010;
		correct = 32'b11101101010100111101110101101010;
		#400 //2.5280273 * -4.098063e+27 = -4.098063e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111000100001000001100101010111;
		b = 32'b01001111101001101101111001100001;
		correct = 32'b01111000100001000001100101010111;
		#400 //2.1434286e+34 * 5599183400.0 = 2.1434286e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111000011100001011010100011;
		b = 32'b10000000011101110111001001010101;
		correct = 32'b01111111000011100001011010100011;
		#400 //1.8886791e+38 * -1.0969439e-38 = 1.8886791e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100011101010000000010100111;
		b = 32'b01011011111011011111101010101011;
		correct = 32'b01011011111011011111101010101011;
		#400 //980.0102 * 1.3397036e+17 = 1.3397036e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101010000100110000110001111;
		b = 32'b10011100000111100000100110010100;
		correct = 32'b00011101000110101101111100101010;
		#400 //2.5726123e-21 * -5.2290194e-22 = 2.0497103e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100100100100111000110000111;
		b = 32'b00110011010010010011101101000110;
		correct = 32'b01001100100100100111000110000111;
		#400 //76778550.0 * 4.685287e-08 = 76778550.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110011011100111100100110111;
		b = 32'b00110101011011000111000111010101;
		correct = 32'b01111110011011100111100100110111;
		#400 //7.924641e+37 * 8.80825e-07 = 7.924641e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101110110100100111110011011;
		b = 32'b11001000011010011100011100000010;
		correct = 32'b11001000011010011100011100000010;
		#400 //-5.778643e-21 * -239388.03 = -239388.03
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001101100101101001011111010;
		b = 32'b11000011000000000001110001100101;
		correct = 32'b11000011000000000001110001100101;
		#400 //-4.3050343e-33 * -128.11092 = -128.11092
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000000011110101101001001001;
		b = 32'b11001011000000010110111101000110;
		correct = 32'b01010000000011110011100111101101;
		#400 //9620235000.0 * -8482630.0 = 9611752000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111101011010111101000100010;
		b = 32'b10100110011000101001010010111111;
		correct = 32'b10110111101011010111101000100010;
		#400 //-2.068008e-05 * -7.861109e-16 = -2.068008e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000011100010100001110000100;
		b = 32'b10000010100111000001110110010000;
		correct = 32'b11010000011100010100001110000100;
		#400 //-16190935000.0 * -2.2939108e-37 = -16190935000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111110101111000010010110010;
		b = 32'b11100011110111110000110001010100;
		correct = 32'b11111111110101111000010010110010;
		#400 //nan * -8.2290245e+21 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011010111000101111010001110;
		b = 32'b00001010101000000110010000011001;
		correct = 32'b01101011010111000101111010001110;
		#400 //2.664102e+26 * 1.5445092e-32 = 2.664102e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111001001111000111000101110;
		b = 32'b00101001110100000111110110011010;
		correct = 32'b00101001110100000111110110011010;
		#400 //1.2605466e-34 * 9.258844e-14 = 9.258844e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001100110111100011000111110;
		b = 32'b01110100110011001100101100111010;
		correct = 32'b11111001100110111001001100001011;
		#400 //-1.0110336e+35 * 1.2980353e+32 = -1.0097355e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101101001000000011011001111;
		b = 32'b01110101000101000110111101111111;
		correct = 32'b01110101000101000110111101111111;
		#400 //1.5424987e-35 * 1.881644e+32 = 1.881644e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011111101001101010010010100;
		b = 32'b00010110000101000100111001010101;
		correct = 32'b11011011111101001101010010010100;
		#400 //-1.3782725e+17 * 1.1980062e-25 = -1.3782725e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010011110111111110111000110;
		b = 32'b11010110001100110011101001001111;
		correct = 32'b11010110001100110011101001001111;
		#400 //-2.2381324e-13 * -49265754000000.0 = -49265754000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001001111000011101110000101;
		b = 32'b11101011011010110001011001011001;
		correct = 32'b11101011011010110001011001011001;
		#400 //2.2657663e-33 * -2.842031e+26 = -2.842031e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011011101110000001101001010;
		b = 32'b01111011110111010100011010001110;
		correct = 32'b01111011010000111000100111010010;
		#400 //-1.282564e+36 * 2.2978572e+36 = 1.0152932e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000111011001111001010111101;
		b = 32'b10111000100000100100100100011001;
		correct = 32'b11010000111011001111001010111101;
		#400 //-31802649000.0 * -6.2124986e-05 = -31802649000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010101000000111111111001111110;
		b = 32'b10100000011111000100101111000001;
		correct = 32'b10100000011111000100101111000011;
		#400 //-2.6655998e-26 * -2.1370295e-19 = -2.1370298e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111100011000010011011110111;
		b = 32'b10100100011001010100001100100110;
		correct = 32'b10100100011001010100001100100110;
		#400 //1.3820075e-29 * -4.9713336e-17 = -4.9713336e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101010110100001011000000110;
		b = 32'b11001111011010100110000010100011;
		correct = 32'b11001111010111001011111101000011;
		#400 //228679780.0 * -3932201700.0 = -3703522000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001110001010011110000100110;
		b = 32'b11101111011110111001000100000111;
		correct = 32'b11101111011110111001000100000111;
		#400 //-4.748259e-33 * -7.7856065e+28 = -7.7856065e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101000111000101101111000111;
		b = 32'b11010100100100011101010110100010;
		correct = 32'b11111101000111000101101111000111;
		#400 //-1.2989756e+37 * -5010835400000.0 = -1.2989756e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010010000010001101110110011001;
		b = 32'b10001110100000001111100000011101;
		correct = 32'b00010010000001111101101110101001;
		#400 //4.3187173e-28 * -3.179336e-30 = 4.286924e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011101011001101011101100000;
		b = 32'b00100000010001110100100110001110;
		correct = 32'b00100000010001111001111111111010;
		#400 //2.8594196e-22 * 1.6880293e-19 = 1.6908887e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100000111110000110111010010;
		b = 32'b11011001110001011111010111001001;
		correct = 32'b11011001110001011111010111001001;
		#400 //0.009707885 * -6965102000000000.0 = -6965102000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110001111000010110001001001;
		b = 32'b11011111111111011101101110001111;
		correct = 32'b11011111111111011101101110001111;
		#400 //-9.961795e-21 * -3.6584743e+19 = -3.6584743e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010011101111010000001011011;
		b = 32'b00010001100001001010010100101001;
		correct = 32'b01100010011101111010000001011011;
		#400 //1.14197515e+21 * 2.0927716e-28 = 1.14197515e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001110110001110110001101110111;
		b = 32'b11101100110110101001000101010111;
		correct = 32'b11101100110110101001000101010111;
		#400 //1672592300.0 * -2.1138574e+27 = -2.1138574e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100111111110111111100111000;
		b = 32'b01100010101001101000111001110111;
		correct = 32'b11111100111111110111111100111000;
		#400 //-1.0612928e+37 * 1.5362126e+21 = -1.0612928e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111101101100010010001000101;
		b = 32'b11000110000110101001011111111011;
		correct = 32'b11010111101101100010010001000101;
		#400 //-400533800000000.0 * -9893.995 = -400533800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011101011101110001001101100;
		b = 32'b01101111101011101011011101111001;
		correct = 32'b01101111101011101011011101111001;
		#400 //-1502246100000.0 * 1.0814439e+29 = 1.0814439e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110101100110111001111010011;
		b = 32'b00000110110110100001010111000101;
		correct = 32'b00100110101100110111001111010011;
		#400 //1.2452014e-15 * 8.2034473e-35 = 1.2452014e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101111011010000111010011001;
		b = 32'b10001010011111100110010110000100;
		correct = 32'b01001101111011010000111010011001;
		#400 //497144600.0 * -1.2248748e-32 = 497144600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101000010100001001001000110;
		b = 32'b00100101110001110000111010110000;
		correct = 32'b01100101000010100001001001000110;
		#400 //4.075148e+22 * 3.453095e-16 = 4.075148e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011001101100011010100000011;
		b = 32'b10011111001100010111110011010010;
		correct = 32'b00110011001101100011010100000011;
		#400 //4.242339e-08 * -3.7584457e-20 = 4.242339e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001010111101010100000110101;
		b = 32'b00111100000101110001010000000100;
		correct = 32'b00111100000101110001010000000100;
		#400 //-4.0895643e-38 * 0.009221081 = 0.009221081
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001110010000011011110110011;
		b = 32'b00001101001011010001111001001101;
		correct = 32'b10110001110010000011011110110011;
		#400 //-5.8270984e-09 * 5.3346214e-31 = -5.8270984e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011000011100010011110100011;
		b = 32'b10010100000110001101010101100011;
		correct = 32'b01001011000011100010011110100011;
		#400 //9316259.0 * -7.716122e-27 = 9316259.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100110101000001101100010001;
		b = 32'b11010101101110011110001010001110;
		correct = 32'b11010101101110011110001010001110;
		#400 //-1.403598e-21 * -25547837000000.0 = -25547837000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000000001011111110100110001;
		b = 32'b11011111001011011001110000011010;
		correct = 32'b11011111001011011001110000011010;
		#400 //-2.0935786 * -1.2509902e+19 = -1.2509902e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001010001011100010100001000;
		b = 32'b01110000101101010000111101011111;
		correct = 32'b01110000101101010000111101011111;
		#400 //12.360603 * 4.4828295e+29 = 4.4828295e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100110001100111000101111010;
		b = 32'b01111000010111001001010000111011;
		correct = 32'b01111000010111001001010000111101;
		#400 //1.9192255e+27 * 1.7895497e+34 = 1.7895499e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000000110010011111010000001;
		b = 32'b11000110100010001111111000100101;
		correct = 32'b11000110100010001111111000100101;
		#400 //-1.2980285e-19 * -17535.072 = -17535.072
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000001111011101101111010110;
		b = 32'b11001000000011001010111011111100;
		correct = 32'b11001000000011001010111011111100;
		#400 //5.7133535e-34 * -144059.94 = -144059.94
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011111100100100000000101010;
		b = 32'b11000111000011001110100001100010;
		correct = 32'b11111011111100100100000000101010;
		#400 //-2.5156745e+36 * -36072.383 = -2.5156745e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110010110001001010011011010;
		b = 32'b01010101111110010011010111001110;
		correct = 32'b01100110010110001001010011011010;
		#400 //2.5569425e+23 * 34251186000000.0 = 2.5569425e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101100010001000011100010110;
		b = 32'b10011011101111001110101010000111;
		correct = 32'b01011101100010001000011100010110;
		#400 //1.229732e+18 * -3.125355e-22 = 1.229732e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101111000111010111100010100000;
		b = 32'b10010010010110011101001110100111;
		correct = 32'b00101111000111010111100010100000;
		#400 //1.4321921e-10 * -6.873401e-28 = 1.4321921e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010100100001001111000110000;
		b = 32'b11101010101010000101101101001001;
		correct = 32'b11101010101010000101101101001001;
		#400 //5.981257e-23 * -1.0176531e+26 = -1.0176531e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000000100101110000110010000;
		b = 32'b11011111001001110011000001001101;
		correct = 32'b11011111001001110011000001001101;
		#400 //5.3435034e-10 * -1.2047214e+19 = -1.2047214e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110011011011001011000101000;
		b = 32'b10101010000111111000011010101101;
		correct = 32'b10101010000111111000011010101101;
		#400 //-1.9192088e-25 * -1.4168762e-13 = -1.4168762e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101110000011011000011110100;
		b = 32'b00011110001010001001111110110101;
		correct = 32'b11001101110000011011000011110100;
		#400 //-406199940.0 * 8.9268726e-21 = -406199940.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100100111101000101010110100;
		b = 32'b01100011100100010111110000000011;
		correct = 32'b11100100011101000101011101100110;
		#400 //-2.3396641e+22 * 5.367428e+21 = -1.8029213e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111110110111100110001000010;
		b = 32'b10111101110110101101010110110110;
		correct = 32'b11011111110110111100110001000010;
		#400 //-3.1676213e+19 * -0.106852934 = -3.1676213e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011011000000111110011000001;
		b = 32'b01110000111000101111110101010010;
		correct = 32'b01110000111000101111110101010010;
		#400 //224.48732 * 5.6199886e+29 = 5.6199886e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001111101000001110000100000;
		b = 32'b10101111100100011000111110001101;
		correct = 32'b10101111100100011000111110001101;
		#400 //2.5240368e-23 * -2.6477345e-10 = -2.6477345e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111100010100010101100001001;
		b = 32'b11001111100001011110111000100011;
		correct = 32'b01011111100010100010101100001001;
		#400 //1.9912123e+19 * -4493952500.0 = 1.9912123e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110001110100110011101000000;
		b = 32'b01000111010110100110011111001111;
		correct = 32'b11010110001110100110011101000000;
		#400 //-51238155000000.0 * 55911.81 = -51238155000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000010110011110101110100101;
		b = 32'b11101110110011100111100101111101;
		correct = 32'b11101110110011100111100101111101;
		#400 //-223150.58 * -3.195039e+28 = -3.195039e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010000001111001010110111111;
		b = 32'b01010000010001110111101011101110;
		correct = 32'b01010000010001110111101011101110;
		#400 //-7.8920825e-09 * 13386889000.0 = 13386889000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011010011101100011110101110;
		b = 32'b11001011101010001011100110011001;
		correct = 32'b11111011010011101100011110101110;
		#400 //-1.0736631e+36 * -22115122.0 = -1.0736631e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100001000000001011111001001;
		b = 32'b11011000101001010011000100100111;
		correct = 32'b11011000101001010011000100100111;
		#400 //3.4714616e-17 * -1453044200000000.0 = -1453044200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010100000011101010010111000;
		b = 32'b10110010100110001000100111000001;
		correct = 32'b10110001001101011010100001001000;
		#400 //1.511431e-08 * -1.7757772e-08 = -2.6434623e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110101000101111101011001011;
		b = 32'b00011001110101100111001100110101;
		correct = 32'b11110110101000101111101011001011;
		#400 //-1.6528101e+33 * 2.2173613e-23 = -1.6528101e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001011001000010111000001100;
		b = 32'b01101001001010011110001110001000;
		correct = 32'b11101000011010010010101000010000;
		#400 //-1.7240784e+25 * 1.2836434e+25 = -4.4043492e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111000011111101110110010111;
		b = 32'b10110010100100111100000011101010;
		correct = 32'b10110010100100111100000011101010;
		#400 //-7.093121e-30 * -1.720078e-08 = -1.720078e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000000001000010100111001000;
		b = 32'b01101011111101110001100001101010;
		correct = 32'b01101011111101110001100001101010;
		#400 //8869323000.0 * 5.9743994e+26 = 5.9743994e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010111100010110110110010111;
		b = 32'b00110111001001111110101101010111;
		correct = 32'b00110111001001111110101101010111;
		#400 //6.5439214e-18 * 1.000877e-05 = 1.000877e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101001101001011100001101101;
		b = 32'b01101100100000000010010101111010;
		correct = 32'b01101101011101001100101100101010;
		#400 //3.4956412e+27 * 1.2393559e+27 = 4.734997e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011111100111101100110001000;
		b = 32'b00100010110110011111101010010100;
		correct = 32'b01100011111100111101100110001000;
		#400 //8.996467e+21 * 5.9083278e-18 = 8.996467e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111010001110101001101000001;
		b = 32'b10111110011101101010001111111111;
		correct = 32'b11101111010001110101001101000001;
		#400 //-6.1688165e+28 * -0.24085997 = -6.1688165e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101010011010001001010110111;
		b = 32'b00011000001110011001110101011111;
		correct = 32'b11101101010011010001001010110111;
		#400 //-3.9666907e+27 * 2.3990142e-24 = -3.9666907e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000001100010001000011100010;
		b = 32'b01001100011011000111100100001100;
		correct = 32'b01100000001100010001000011100010;
		#400 //5.1035785e+19 * 61989936.0 = 5.1035785e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011001000110110001100000001;
		b = 32'b00000110110000001011101011000110;
		correct = 32'b00111011001000110110001100000001;
		#400 //0.0024930837 * 7.249681e-35 = 0.0024930837
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101111000111111011101000001;
		b = 32'b10100100101100100110001101100010;
		correct = 32'b11001101111000111111011101000001;
		#400 //-478079000.0 * -7.7363556e-17 = -478079000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000101010111010000001001000;
		b = 32'b10010010010010110101110111101100;
		correct = 32'b11101000101010111010000001001000;
		#400 //-6.4838507e+24 * -6.4171273e-28 = -6.4838507e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000101010011100011001100100;
		b = 32'b01110000001110010100000101011010;
		correct = 32'b11110000000110100100101101101110;
		#400 //-4.2034245e+29 * 2.2933493e+29 = -1.9100752e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001110011000010100100011100;
		b = 32'b00100000000000000110111001100000;
		correct = 32'b00100000000000000110111001100000;
		#400 //-7.4996754e-38 * 1.0878542e-19 = 1.0878542e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110110011101011110011010100;
		b = 32'b10011010101010101001000011110001;
		correct = 32'b00100110110011101011110011010011;
		#400 //1.4345303e-15 * -7.054452e-23 = 1.4345302e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001111010010000011110011010;
		b = 32'b01110000010110111100001011000110;
		correct = 32'b01111001111010010000011110110101;
		#400 //1.5124492e+35 * 2.7205074e+29 = 1.5124519e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101111010000011111011101100;
		b = 32'b00101001001111001111101100001001;
		correct = 32'b00101001001111001111101100001011;
		#400 //6.147495e-21 * 4.1962124e-14 = 4.196213e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001110011110010001011000001110;
		b = 32'b11001110000110011101000010110001;
		correct = 32'b01001101101111101000101010111010;
		#400 //1044743040.0 * -645147700.0 = 399595330.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000000100100101001100100100;
		b = 32'b11011000000010000101011111101001;
		correct = 32'b11011000000010000101011111101001;
		#400 //4.403301e-34 * -599644600000000.0 = -599644600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010100110010001010010010111;
		b = 32'b10111101111110000010010111111000;
		correct = 32'b10111101111110000010010111111000;
		#400 //6.331258e-23 * -0.12116617 = -0.12116617
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001110000111010011001011010010;
		b = 32'b00110100110010100101101010110111;
		correct = 32'b00110100110010100101101010110111;
		#400 //1.9376213e-30 * 3.7691436e-07 = 3.7691436e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111001101000010101010101111;
		b = 32'b00110100101110111110111100110001;
		correct = 32'b00110100101110111110111100110001;
		#400 //1.3554239e-34 * 3.50055e-07 = 3.50055e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000000111111001010100010011;
		b = 32'b00100011000000001100000111101011;
		correct = 32'b00100011000000110100000000111111;
		#400 //1.3517148e-19 * 6.979958e-18 = 7.115129e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010000011110101111000100000;
		b = 32'b00000010011100110100101010110100;
		correct = 32'b00001010000011110101111100010011;
		#400 //6.9029025e-33 * 1.7874259e-37 = 6.903081e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110101111011011000111001010;
		b = 32'b00101011000110010011001011011111;
		correct = 32'b11001110101111011011000111001010;
		#400 //-1591272700.0 * 5.4427117e-13 = -1591272700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101010101100100010011001110;
		b = 32'b10000111100001111110010110001011;
		correct = 32'b11001101010101100100010011001110;
		#400 //-224677090.0 * -2.0447456e-34 = -224677090.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111010100101111010111011111;
		b = 32'b11011000010001010111111000010000;
		correct = 32'b11011000010001010111111000010000;
		#400 //54005.87 * -868580900000000.0 = -868580900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101111110101011000110101001101;
		b = 32'b11111100011001000001101000011101;
		correct = 32'b11111100011001000001101000011101;
		#400 //3.8844875e-10 * -4.7374933e+36 = -4.7374933e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000111011100100100100111110;
		b = 32'b01010110010101001011010110101011;
		correct = 32'b01100000111011100100100101000101;
		#400 //1.3736259e+20 * 58469180000000.0 = 1.3736265e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010011000000100100000100001;
		b = 32'b00010100010001011111111000101010;
		correct = 32'b10101010011000000100100000100001;
		#400 //-1.9920221e-13 * 9.996083e-27 = -1.9920221e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010010000110010000001011100;
		b = 32'b10001100000101000111101010000010;
		correct = 32'b11001010010000110010000001011100;
		#400 //-3196951.0 * -1.1438371e-31 = -3196951.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000000010000000001110111001;
		b = 32'b10100111010110101100111111111001;
		correct = 32'b10100111010110101100111111111001;
		#400 //-7.3602e-40 * -3.036632e-15 = -3.036632e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001000000110111101110101001;
		b = 32'b00011011011010110111001010110111;
		correct = 32'b11001001000000110111101110101001;
		#400 //-538554.56 * 1.9475811e-22 = -538554.56
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100101111110001010011110101;
		b = 32'b01001101010010110110000101110011;
		correct = 32'b01001101010010110110000101110011;
		#400 //8.286855e-17 * 213260080.0 = 213260080.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010110100000001010100011000;
		b = 32'b01001011010010000101110011011100;
		correct = 32'b01001011010010000101110011011100;
		#400 //-2.422398e-08 * 13130972.0 = 13130972.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110010101001101101110111101;
		b = 32'b11010111001110000000011010110001;
		correct = 32'b11100110010101001101101110111101;
		#400 //-2.5129879e+23 * -202338880000000.0 = -2.5129879e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100111101000011011001010101;
		b = 32'b00100100010001000101101000110100;
		correct = 32'b00110100111101000011011001010101;
		#400 //4.5488073e-07 * 4.257713e-17 = 4.5488073e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000011100000101001100111110;
		b = 32'b00001001110100110010001101101000;
		correct = 32'b11000000011100000101001100111110;
		#400 //-3.7550807 * 5.0829698e-33 = -3.7550807
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010110000011110100110100001;
		b = 32'b01111100101101111111100111001011;
		correct = 32'b01111100101101111111100111001011;
		#400 //-8.020038e-23 * 7.642054e+36 = 7.642054e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010111101100110000101010010;
		b = 32'b00110011000110000110010011101011;
		correct = 32'b01001010111101100110000101010010;
		#400 //8073385.0 * 3.5482042e-08 = 8073385.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000010000100100110100011010;
		b = 32'b01100111110001110100010011011011;
		correct = 32'b01100111110001110100010011011011;
		#400 //-198964.4 * 1.8820422e+24 = 1.8820422e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100001101010100011000110011;
		b = 32'b11100000101001100100101010111101;
		correct = 32'b11100000101001100100101010111101;
		#400 //3.930758e-17 * -9.586078e+19 = -9.586078e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010101111101110001001101000;
		b = 32'b01110111011100011110011010010011;
		correct = 32'b01110111011100011110011010010011;
		#400 //-6254900.0 * 4.9063287e+33 = 4.9063287e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111100111100101101000011001;
		b = 32'b01100111101011101001010101100100;
		correct = 32'b01100111101011101001010101100100;
		#400 //81076.195 * 1.6488951e+24 = 1.6488951e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100100110101011101110100001001;
		b = 32'b11010100100011000001100011000001;
		correct = 32'b11010100100011000001100011000001;
		#400 //-9.274847e-17 * -4813686000000.0 = -4813686000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011010000101010101010101000;
		b = 32'b10000010001000010000100100100011;
		correct = 32'b00100011010000101010101010101000;
		#400 //1.0552899e-17 * -1.1831034e-37 = 1.0552899e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000001010011110111110100000;
		b = 32'b11010011001101110011011110110101;
		correct = 32'b11010011001110011101111101110100;
		#400 //-11404214000.0 * -786913600000.0 = -798317900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000011000111011111010110100;
		b = 32'b11011001100000010011100101100101;
		correct = 32'b11011001100000010011100101100101;
		#400 //-5.4298624e-05 * -4546672000000000.0 = -4546672000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010011010001111010111111001;
		b = 32'b10100101111010111110111000110011;
		correct = 32'b01011010011010001111010111111001;
		#400 //1.6393161e+16 * -4.0927412e-16 = 1.6393161e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101110011111001110101010000;
		b = 32'b10001000000110011000110001111110;
		correct = 32'b11100101110011111001110101010000;
		#400 //-1.2255397e+23 * -4.620691e-34 = -1.2255397e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011100010111000000000010000;
		b = 32'b11000111011100001011110100011110;
		correct = 32'b11000111011100001011110100011110;
		#400 //2.307838e-22 * -61629.117 = -61629.117
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010011110001010110001011101;
		b = 32'b00001010111011011110001111110001;
		correct = 32'b11110010011110001010110001011101;
		#400 //-4.925482e+30 * 2.2908012e-32 = -4.925482e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101010011110110101100000001;
		b = 32'b01100011111111101111010001111100;
		correct = 32'b01100011111111101111010001111100;
		#400 //-7.726922e-07 * 9.40618e+21 = 9.40618e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111001101010100010011101000;
		b = 32'b01000100000111000110101111000111;
		correct = 32'b01000100000111000011111001110110;
		#400 //-0.7080827 * 625.684 = 624.97595
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101101001001111100001011110;
		b = 32'b01010100100101001110100011111101;
		correct = 32'b11010101011111110111110000111110;
		#400 //-22673330000000.0 * 5116512400000.0 = -17556818000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001010010001101101101010010;
		b = 32'b10000111111101101001010101010010;
		correct = 32'b00001001001010100000100010101000;
		#400 //2.4177248e-33 * -3.7101729e-34 = 2.0467076e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000100111111000100111011111;
		b = 32'b01110111011011000010101111011110;
		correct = 32'b01110111011011000010101111011110;
		#400 //4.98558 * 4.7901242e+33 = 4.7901242e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011101000001100100010101111;
		b = 32'b10000000111010111101010100011110;
		correct = 32'b10101011101000001100100010101111;
		#400 //-1.1424385e-12 * -2.1657794e-38 = -1.1424385e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111100100001110111111001100;
		b = 32'b11100011000111000010101010111100;
		correct = 32'b11100011000111000010101010111100;
		#400 //-4863269000.0 * -2.8807714e+21 = -2.8807714e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111000001010010010100010010100;
		b = 32'b01101011101101111010001100110000;
		correct = 32'b01111000001010010010100010010100;
		#400 //1.3723769e+34 * 4.440081e+26 = 1.3723769e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010010101110011010000010001;
		b = 32'b01100000111000011000100111101100;
		correct = 32'b01110010010101110011010000010001;
		#400 //4.2625422e+30 * 1.3001424e+20 = 4.2625422e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110110001000010001110100101;
		b = 32'b11001011011111000010000111011101;
		correct = 32'b11001011011111000010000111011101;
		#400 //-1.3609894e-15 * -16523741.0 = -16523741.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111111101111010110001111001;
		b = 32'b11100011110010110011100101111001;
		correct = 32'b11100011110010110011100101111001;
		#400 //1.6005539e-24 * -7.497661e+21 = -7.497661e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010110000011001000001100001;
		b = 32'b11001101000010100100100010100100;
		correct = 32'b11110010110000011001000001100001;
		#400 //-7.667859e+30 * -145001020.0 = -7.667859e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111010011111011000001100010000;
		b = 32'b11100100100010000011011100110011;
		correct = 32'b11100100100010000011011100110011;
		#400 //0.0009670714 * -2.0101878e+22 = -2.0101878e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011010110111110100000011001;
		b = 32'b10001101001110111011010100111001;
		correct = 32'b00110011010110111110100000011001;
		#400 //5.1201003e-08 * -5.7841963e-31 = 5.1201003e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100000101010111110011011100;
		b = 32'b11100001111111100011010110111111;
		correct = 32'b01100100000011011000101100101110;
		#400 //1.1030248e+22 * -5.8616823e+20 = 1.044408e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111011100100111111111101110;
		b = 32'b10011100111000010110110001000011;
		correct = 32'b01000111011100100111111111101110;
		#400 //62079.93 * -1.4917236e-21 = 62079.93
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111100100111010111111000111;
		b = 32'b00101000110101001011011110111101;
		correct = 32'b00101000111110011010001110101111;
		#400 //4.0991274e-15 * 2.3616412e-14 = 2.771554e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110101100010011000011101001;
		b = 32'b01001001111101010011000101101101;
		correct = 32'b01001001111101010011000101101101;
		#400 //-1.2295099e-15 * 2008621.6 = 2008621.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000111110101110111010000001;
		b = 32'b00101101010110101100001110100100;
		correct = 32'b11011000111110101110111010000001;
		#400 //-2207218200000000.0 * 1.2435306e-11 = -2207218200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001000001111101000100000001100;
		b = 32'b10001001100001001011000000101111;
		correct = 32'b10001001100111001000000100110000;
		#400 //-5.7335968e-34 * -3.1943526e-33 = -3.767712e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011111010011110001110100110;
		b = 32'b11111011010011110000100010000111;
		correct = 32'b11111011010011110000100010000111;
		#400 //-30656332.0 * -1.0749784e+36 = -1.0749784e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111010100010101100010001000;
		b = 32'b11010110100010011001011011110000;
		correct = 32'b11010110100010011001010101001101;
		#400 //3512240000.0 * -75640680000000.0 = -75637170000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011100010100001010010011001110;
		b = 32'b01010001001101100011110100010010;
		correct = 32'b01010001001101100011110100010010;
		#400 //6.903443e-22 * 48919290000.0 = 48919290000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101100101001011110110101100110;
		b = 32'b01001010010010011100100100110001;
		correct = 32'b01001010010010011100100100110001;
		#400 //4.7159386e-12 * 3306060.2 = 3306060.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001101000101111111000001010;
		b = 32'b01100100000111010010000111110110;
		correct = 32'b01100100000111010010000111110110;
		#400 //20.374043 * 1.1594344e+22 = 1.1594344e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010110110010001010111001000;
		b = 32'b00011001000111011100011101001001;
		correct = 32'b11000010110110010001010111001000;
		#400 //-108.54254 * 8.156955e-24 = -108.54254
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110010010001001011000011110;
		b = 32'b00011101101000010000010110001010;
		correct = 32'b01010110010010001001011000011110;
		#400 //55136770000000.0 * 4.2622072e-21 = 55136770000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111000010111100011101000000;
		b = 32'b11110001110001001100101000010011;
		correct = 32'b11110001110001001100101000010011;
		#400 //-2345091000.0 * -1.9489073e+30 = -1.9489073e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010111010001001101000100001;
		b = 32'b00011001100111011010010010100101;
		correct = 32'b00011001100111011010010010100101;
		#400 //3.4177802e-37 * 1.6299919e-23 = 1.6299919e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111010111001111110100011111;
		b = 32'b10011001110110111100011110111111;
		correct = 32'b10011001110110111100011111000110;
		#400 //-1.0895587e-29 * -2.2724746e-23 = -2.2724757e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011110010000101101001011110;
		b = 32'b00100010101111111101001000011101;
		correct = 32'b00100010101111111100111011111100;
		#400 //-3.3145623e-22 * 5.199312e-18 = 5.1989807e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101101011110010111000111110;
		b = 32'b11110001010100011111010100101110;
		correct = 32'b11110001010100011111010100101110;
		#400 //4.6369928e-21 * -1.0396603e+30 = -1.0396603e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100101010100111001001001101;
		b = 32'b00101001110101011101111100111011;
		correct = 32'b00110100101010100111001001010000;
		#400 //3.1748132e-07 * 9.4978245e-14 = 3.174814e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000101001011000011111101001;
		b = 32'b11010001111101000111011110101110;
		correct = 32'b11010001111101000111011110101110;
		#400 //6.529043e-29 * -131247490000.0 = -131247490000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100000101100010100100010010;
		b = 32'b00100001110100100110101110001111;
		correct = 32'b00100001110100100110101110001111;
		#400 //-7.581164e-27 * 1.4258624e-18 = 1.4258624e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110010010111010101100100100;
		b = 32'b10011111010101000101000110010101;
		correct = 32'b10100110010010111010111001110101;
		#400 //-7.066171e-16 * -4.496023e-20 = -7.0666206e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001010111100111001010100110;
		b = 32'b00001110100011010010110110101100;
		correct = 32'b01010001010111100111001010100110;
		#400 //59712890000.0 * 3.4803164e-30 = 59712890000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001011011001011010100101001;
		b = 32'b01101111001011010010000100011000;
		correct = 32'b01101111001011010010000100011000;
		#400 //3.4445498e-09 * 5.3580915e+28 = 5.3580915e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000011110000110110001011100;
		b = 32'b10010101000011111000011001111101;
		correct = 32'b10111000011110000110110001011100;
		#400 //-5.9228725e-05 * -2.8984713e-26 = -5.9228725e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011011111000001111011011001;
		b = 32'b10100111111111110111110110010111;
		correct = 32'b10100111111111110111110110010111;
		#400 //2.0854919e-22 * -7.0912883e-15 = -7.0912883e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011010000011000000100100011;
		b = 32'b10110010100101111010100111111011;
		correct = 32'b01011011010000011000000100100011;
		#400 //5.4466658e+16 * -1.7656012e-08 = 5.4466658e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111111001001010001100110000;
		b = 32'b00111010011101110110011110011001;
		correct = 32'b00111010011101110110011110011001;
		#400 //1.4775349e-24 * 0.00094377395 = 0.00094377395
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101100110101001011011010011;
		b = 32'b01100111000010100001000100111100;
		correct = 32'b01110101100110101001011011010011;
		#400 //3.9193008e+32 * 6.520045e+23 = 3.9193008e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000110110100111100010010000;
		b = 32'b10001110111011110010001100001111;
		correct = 32'b11110000110110100111100010010000;
		#400 //-5.4090787e+29 * -5.895181e-30 = -5.4090787e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111000010010110010001111101;
		b = 32'b10101000110001100010111110101011;
		correct = 32'b11010111000010010110010001111101;
		#400 //-151064690000000.0 * -2.2003089e-14 = -151064690000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000110000000111010111011001101;
		b = 32'b01001100110111010101100011100111;
		correct = 32'b01001100110111010101100011100111;
		#400 //-2.4766785e-35 * 116049720.0 = 116049720.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101100001101110011011100011;
		b = 32'b00110111110100110100011110010111;
		correct = 32'b01001101100001101110011011100011;
		#400 //282909800.0 * 2.5186497e-05 = 282909800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111100010110111111000100100;
		b = 32'b00011111110101000100101101100100;
		correct = 32'b01100111100010110111111000100100;
		#400 //1.3174716e+24 * 8.9910216e-20 = 1.3174716e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110001001111101011011100011;
		b = 32'b11111001111011111011011001011111;
		correct = 32'b11111001111011111011011001011111;
		#400 //-703969500.0 * -1.5558223e+35 = -1.5558223e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001010110000000000111010011;
		b = 32'b00001011001011100100011000101100;
		correct = 32'b01000001010110000000000111010011;
		#400 //13.500445 * 3.3563972e-32 = 13.500445
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011111101010010011000111110;
		b = 32'b10111110110111000010100100110111;
		correct = 32'b01101011111101010010011000111110;
		#400 //5.9273484e+26 * -0.43000194 = 5.9273484e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111110100111010010111110100;
		b = 32'b11100100010000010110001110100101;
		correct = 32'b11100100010000010110001110100101;
		#400 //1.3677448e-24 * -1.4269607e+22 = -1.4269607e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000001101011000111111101110;
		b = 32'b00110101001000101100000011001011;
		correct = 32'b10111000001100110000010011101011;
		#400 //-4.3287808e-05 * 6.0630254e-07 = -4.2681506e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011000000010011111111111111;
		b = 32'b00110101100010110001001100100001;
		correct = 32'b00110101100010110001001100100001;
		#400 //1.6313642e-27 * 1.0361874e-06 = 1.0361874e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101000010100001001000100000;
		b = 32'b10101011111100010011101011001100;
		correct = 32'b10111101000010100001001000100000;
		#400 //-0.03370869 * -1.7140399e-12 = -0.03370869
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001010001010111010011101111;
		b = 32'b11101101011010110110101111111101;
		correct = 32'b11101101011010110110101111111101;
		#400 //6.6900957e-19 * -4.5537204e+27 = -4.5537204e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111010001100011101001101001;
		b = 32'b01100010010000100000010000010010;
		correct = 32'b01100010010000100000010000010010;
		#400 //1.1815319e-05 * 8.947404e+20 = 8.947404e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100010010001010101110110000001;
		b = 32'b00001000100001101100111100101001;
		correct = 32'b11100010010001010101110110000001;
		#400 //-9.1018656e+20 * 8.113535e-34 = -9.1018656e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010110000001111111001111101;
		b = 32'b11001100011101001011111110010101;
		correct = 32'b01011010110000001111111001111101;
		#400 //2.7161504e+16 * -64159316.0 = 2.7161504e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010111100100010111101000111;
		b = 32'b10000001111010111110100111010000;
		correct = 32'b10001010111100100010111110000010;
		#400 //-2.3321536e-32 * -8.666087e-38 = -2.3321623e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110001110001101001010011100;
		b = 32'b10101111011110000111010010011101;
		correct = 32'b10111110001110001101001010011100;
		#400 //-0.18049091 * -2.2596898e-10 = -0.18049091
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111010001001010000100100110;
		b = 32'b11010100101011001110001010011000;
		correct = 32'b11010100101011001110001010011000;
		#400 //-0.76808393 * -5940288000000.0 = -5940288000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000110000111011111100101101;
		b = 32'b00110110001101110000111110010000;
		correct = 32'b00110110001101110000111110010000;
		#400 //-3.3160794e-19 * 2.7278184e-06 = 2.7278184e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110010001010111100101111001;
		b = 32'b00000011100000011011110000010010;
		correct = 32'b10110110010001010111100101111001;
		#400 //-2.9425994e-06 * 7.625117e-37 = -2.9425994e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101010010011000011110010000011;
		b = 32'b01110011100010001100110010011000;
		correct = 32'b01110011100010001100110010011000;
		#400 //1.8139834e-13 * 2.1676698e+31 = 2.1676698e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001111011111010110000000110;
		b = 32'b10110011010111111000101101000001;
		correct = 32'b10110011010111111000101101000001;
		#400 //5.7698927e-33 * -5.2047884e-08 = -5.2047884e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001110110101110101010000110;
		b = 32'b10001101000111111000110110010001;
		correct = 32'b11111001110110101110101010000110;
		#400 //-1.4208468e+35 * -4.916606e-31 = -1.4208468e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101000111011100101111000101000;
		b = 32'b00111001101100001000110110001111;
		correct = 32'b00111001101100001000110110001111;
		#400 //2.6464142e-14 * 0.00033674805 = 0.00033674805
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001001110011011011100101010;
		b = 32'b00011111001011101110001100011010;
		correct = 32'b01111001001110011011011100101010;
		#400 //6.026812e+34 * 3.7033787e-20 = 6.026812e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010110001111111110010111111;
		b = 32'b10001001011011000001001110100110;
		correct = 32'b01110010110001111111110010111111;
		#400 //7.922313e+30 * -2.8416705e-33 = 7.922313e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011001001111111010010111001111;
		b = 32'b00101000101100000100001110001010;
		correct = 32'b00101000101100000100001110001010;
		#400 //-9.907953e-24 * 1.9569216e-14 = 1.9569216e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101011100101110011111001010;
		b = 32'b11010010100000110100000000110000;
		correct = 32'b01010101011011101100110111001000;
		#400 //16692334000000.0 * -281858800000.0 = 16410474000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110000011101100110010010111;
		b = 32'b10101010101111010111111011100110;
		correct = 32'b01010110000011101100110010010111;
		#400 //39252340000000.0 * -3.3661198e-13 = 39252340000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000101100110001001000011011;
		b = 32'b01010100111000101011111100100000;
		correct = 32'b01010100111000101011111100100001;
		#400 //366736.84 * 7790953000000.0 = 7790954000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011100100011011101011111000;
		b = 32'b01010000111111101101001011001111;
		correct = 32'b01010000111111101101001011001111;
		#400 //-3.678751e-27 * 34201827000.0 = 34201827000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101001110011110000001011111;
		b = 32'b10000100011000001000100111011010;
		correct = 32'b01100101001110011110000001011111;
		#400 //5.4861045e+22 * -2.6394372e-36 = 5.4861045e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111101111000010000101010101;
		b = 32'b01010110100000100001000111110010;
		correct = 32'b01010110100000100001000111110010;
		#400 //96322.664 * 71506790000000.0 = 71506790000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011001011011111100110111100;
		b = 32'b01111100001011010001110000101011;
		correct = 32'b01111100001011010001110000101011;
		#400 //-2.103235e+26 * 3.5953547e+36 = 3.5953547e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110111100011100001010111010;
		b = 32'b11100100110010100101010111001110;
		correct = 32'b11100100110010100110010011101010;
		#400 //-8.7103454e+18 * -2.9859401e+22 = -2.9868111e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110000100100000111010001010;
		b = 32'b10010100011111011111111000011001;
		correct = 32'b11001110000100100000111010001010;
		#400 //-612606600.0 * -1.2823348e-26 = -612606600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010110011111101001100101111;
		b = 32'b01010110011010111011110000101001;
		correct = 32'b01010110011010111011110000101001;
		#400 //3.053713e-37 * 64798344000000.0 = 64798344000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010100100010001111001011001;
		b = 32'b01100110100101111000010101001011;
		correct = 32'b01100110100101111000010101001011;
		#400 //-3.933446e-18 * 3.5776808e+23 = 3.5776808e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010101000101001010001001110;
		b = 32'b11111000000000101110100110010011;
		correct = 32'b11111000000000101110100110010011;
		#400 //4.406721e-18 * -1.0620876e+34 = -1.0620876e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101001101010110110100111110;
		b = 32'b01011010100001010100111011110011;
		correct = 32'b01011010100001010100111011110011;
		#400 //-2.4011627e-21 * 1.8761489e+16 = 1.8761489e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000010100110001000000001011;
		b = 32'b11010000000011110111110001011111;
		correct = 32'b11010000000011110111110001011111;
		#400 //-2.727921e-24 * -9629171000.0 = -9629171000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010101100110000010111011111;
		b = 32'b10101011001111111010110011111101;
		correct = 32'b11000010101100110000010111011111;
		#400 //-89.51147 * -6.80969e-13 = -89.51147
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011100110100110011110001010;
		b = 32'b10000100011010111000110000000110;
		correct = 32'b10101011100110100110011110001010;
		#400 //-1.0971096e-12 * -2.7688413e-36 = -1.0971096e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101111001000001000111110000;
		b = 32'b00111110101000010110110010111101;
		correct = 32'b00111110101000010110110010111101;
		#400 //-3.956385e-16 * 0.31528273 = 0.31528273
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011110101011110001111010110;
		b = 32'b00101100100100011100111010100011;
		correct = 32'b11001011110101011110001111010110;
		#400 //-28034988.0 * 4.144089e-12 = -28034988.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111010110010011000010100000;
		b = 32'b11110011110101000010100011001011;
		correct = 32'b11110011110101000010100011001011;
		#400 //7.0177855e-25 * -3.361799e+31 = -3.361799e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111001110100001000001000101;
		b = 32'b11101001000011001101011001001001;
		correct = 32'b01111111001110100001000001000101;
		#400 //2.4732088e+38 * -1.0641347e+25 = 2.4732088e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001000000101011111110000000;
		b = 32'b01101000010101111100110011110101;
		correct = 32'b01101000010101111100110011110101;
		#400 //2300144000000000.0 * 4.0763583e+24 = 4.0763583e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000100011010001001000010111;
		b = 32'b11111000000100110100010010100100;
		correct = 32'b11111000000100110100010010100100;
		#400 //-5.5642566e-29 * -1.194781e+34 = -1.194781e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011110111001110010010010101;
		b = 32'b00000101110000010011101010001101;
		correct = 32'b01011011110111001110010010010101;
		#400 //1.2435165e+17 * 1.8171141e-35 = 1.2435165e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000000000001100001010100100;
		b = 32'b00010000010101111101111011111101;
		correct = 32'b10011000000000001100000111001100;
		#400 //-1.664188e-24 * 4.2573058e-29 = -1.6641455e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100000001101101111100110011;
		b = 32'b10110110100010011111000010010110;
		correct = 32'b10110110100010011111000010010110;
		#400 //1.0390151e-31 * -4.110926e-06 = -4.110926e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110000001001110111110101001;
		b = 32'b01010100010101111000111110001001;
		correct = 32'b01010100010101111000111110001001;
		#400 //2.5002515e-35 * 3703304400000.0 = 3703304400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010011101101100111110011001101;
		b = 32'b01110011000011010000110001110111;
		correct = 32'b01110011000011010000110001110111;
		#400 //1567555700000.0 * 1.1175029e+31 = 1.1175029e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110101010001001010111111000;
		b = 32'b00000101101100111101101110011001;
		correct = 32'b11000110101010001001010111111000;
		#400 //-21578.984 * 1.6913747e-35 = -21578.984
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000010111011000001100110001;
		b = 32'b10001001110000001110111110000011;
		correct = 32'b10111000010111011000001100110001;
		#400 //-5.2812687e-05 * -4.6447554e-33 = -5.2812687e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010010110011111010110011010001;
		b = 32'b10000001101111000000100111001101;
		correct = 32'b00010010110011111010110011010001;
		#400 //1.3106139e-27 * -6.9074357e-38 = 1.3106139e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100110110011111111101011001;
		b = 32'b11011011011010100101110001101000;
		correct = 32'b11111100110110011111111101011001;
		#400 //-9.05526e+36 * -6.5966746e+16 = -9.05526e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110001001000011001101000100;
		b = 32'b11000010000110101011001110000001;
		correct = 32'b11000010000110101011001110000001;
		#400 //-5.696841e-16 * -38.675297 = -38.675297
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101001001111010101100011100;
		b = 32'b11111111111101001010010011110101;
		correct = 32'b11111111111101001010010011110101;
		#400 //1.4542915e-16 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101010110111000100111101000;
		b = 32'b11011110011100010011100111000101;
		correct = 32'b11101101010110111000100111101000;
		#400 //-4.246496e+27 * -4.3455352e+18 = -4.246496e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100001101000111100011111100;
		b = 32'b10111110000110101110000101000110;
		correct = 32'b11010100001101000111100011111100;
		#400 //-3100495600000.0 * -0.15124997 = -3100495600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111101001001010110111111110;
		b = 32'b00000010111011100111011010001101;
		correct = 32'b11101111101001001010110111111110;
		#400 //-1.0193177e+29 * 3.5039002e-37 = -1.0193177e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110110001101100000000011011;
		b = 32'b01101000010111110101000110011011;
		correct = 32'b01101000010111110101000110011011;
		#400 //109264195000000.0 * 4.2183723e+24 = 4.2183723e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101001100101110110001100000;
		b = 32'b10100111111100110110000000111100;
		correct = 32'b00111101001100101110110001100000;
		#400 //0.043682456 * -6.7550386e-15 = 0.043682456
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010100001011000010011101000;
		b = 32'b01110111110101011100100001001011;
		correct = 32'b01110111110101011110100110101100;
		#400 //5.289239e+30 * 8.672044e+33 = 8.677333e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101110100011010011110111110;
		b = 32'b10001111101011111011100100010000;
		correct = 32'b01111101110100011010011110111110;
		#400 //3.4834952e+37 * -1.7327616e-29 = 3.4834952e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110111101010111100001001001;
		b = 32'b11010110111111101000011100101000;
		correct = 32'b11110110111101010111100001001001;
		#400 //-2.4893602e+33 * -139928220000000.0 = -2.4893602e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001111111110100001010110001;
		b = 32'b10110011101001001011111110111110;
		correct = 32'b01011001111111110100001010110001;
		#400 //8981181000000000.0 * -7.671723e-08 = 8981181000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001111011001011100001001100;
		b = 32'b01001000110001010100000101011111;
		correct = 32'b11010001111011001011100000011011;
		#400 //-127088030000.0 * 403978.97 = -127087630000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101000001111111111110010010001;
		b = 32'b11100011001101111000011011110001;
		correct = 32'b11100011001101111000011011110001;
		#400 //1.06573965e-14 * -3.3854777e+21 = -3.3854777e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011001110110001001010111010;
		b = 32'b10000010110011011110110010010110;
		correct = 32'b00001011001110110001001001010011;
		#400 //3.6028978e-32 * -3.0257836e-37 = 3.6028676e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010100101001100100010010100;
		b = 32'b10000101101111000101000010100010;
		correct = 32'b01111010100101001100100010010100;
		#400 //3.8626407e+35 * -1.7709055e-35 = 3.8626407e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100011011100010010111001101101;
		b = 32'b11111000011011001101010111000000;
		correct = 32'b11111000011011001101010111000000;
		#400 //-1.3074467e-17 * -1.9214335e+34 = -1.9214335e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101101010011101000110011110;
		b = 32'b10011011100100110001111100100011;
		correct = 32'b10011011100100110001111100100011;
		#400 //-1.5969685e-35 * -2.4339232e-22 = -2.4339232e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101000001101101110111110011;
		b = 32'b00000111101001110000000011101010;
		correct = 32'b11101101000001101101110111110011;
		#400 //-2.608707e+27 * 2.5127904e-34 = -2.608707e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100100010110100111111000010010;
		b = 32'b00100010011111110100010101010011;
		correct = 32'b10100100010010101000100110111101;
		#400 //-4.7378e-17 * 3.4595644e-18 = -4.3918437e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011111011111110100101001100;
		b = 32'b10100101110011011111011111001100;
		correct = 32'b10110011111011111110100101001100;
		#400 //-1.1171741e-07 * -3.5729745e-16 = -1.1171741e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011101111001101111001001000;
		b = 32'b01110001001000001010101111101110;
		correct = 32'b01110001001000001010101111101110;
		#400 //-4.767706e-27 * 7.956072e+29 = 7.956072e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001111111110100000010110010;
		b = 32'b00101111010001111010110001110100;
		correct = 32'b01000001111111110100000010110010;
		#400 //31.90659 * 1.8160212e-10 = 31.90659
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100100010101111000001011010;
		b = 32'b11010110011100111101000111100010;
		correct = 32'b11110100100010101111000001011010;
		#400 //-8.806297e+31 * -67020690000000.0 = -8.806297e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011011011001110011000110000;
		b = 32'b11101100000111000110011000100001;
		correct = 32'b11101100000111000110011000100001;
		#400 //2.9900879e-27 * -7.562989e+26 = -7.562989e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111111011110001010101000111;
		b = 32'b11100101011111101011010110011000;
		correct = 32'b11100101011111101011010110011000;
		#400 //-525749330000000.0 * -7.517693e+22 = -7.517693e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000101110010100110100000010;
		b = 32'b00011010010101001010001001110100;
		correct = 32'b01010000101110010100110100000010;
		#400 //24870654000.0 * 4.39718e-23 = 24870654000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001011110000111000011100000;
		b = 32'b10100110111010101100001111110001;
		correct = 32'b01001001011110000111000011100000;
		#400 //1017614.0 * -1.6290122e-15 = 1017614.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101000010110100001011110000;
		b = 32'b01011100000100100111101011111011;
		correct = 32'b01011101001011111110000110101111;
		#400 //6.271779e+17 * 1.6492226e+17 = 7.921002e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011101001100110101000000010;
		b = 32'b01110001010010000011011101000010;
		correct = 32'b01110001010010000011011101000010;
		#400 //-2.7530902e-22 * 9.914209e+29 = 9.914209e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111000100101100000110011010;
		b = 32'b00000000010001110011011011100001;
		correct = 32'b11101111000100101100000110011010;
		#400 //-4.541886e+28 * 6.540007e-39 = -4.541886e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001011011111011100010110101;
		b = 32'b01000111100001110001100100100011;
		correct = 32'b01001001100000000100110111101101;
		#400 //981899.3 * 69170.27 = 1051069.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000010000101000001000011100;
		b = 32'b10110011100010111000110100101000;
		correct = 32'b01110000010000101000001000011100;
		#400 //2.4078954e+29 * -6.498368e-08 = 2.4078954e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011111011101101010100001100;
		b = 32'b01101000000111001110110011110100;
		correct = 32'b01101000000111001110110011110100;
		#400 //3.9511475e-22 * 2.9642407e+24 = 2.9642407e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101010011001010111000010111;
		b = 32'b10111010110001101001101110110010;
		correct = 32'b01101101010011001010111000010111;
		#400 //3.9590877e+27 * -0.0015152602 = 3.9590877e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010111010100000101001101011111;
		b = 32'b11010001100001001100101110110101;
		correct = 32'b11010001100001001100101110110101;
		#400 //-6.7313654e-25 * -71294165000.0 = -71294165000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111010000111111000100010100;
		b = 32'b00001111001100011100101010101101;
		correct = 32'b01010111010000111111000100010100;
		#400 //215440190000000.0 * 8.765808e-30 = 215440190000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110111001011101111001011111;
		b = 32'b11100100111001110100001110010011;
		correct = 32'b11101110111001011101111001101101;
		#400 //-3.5570449e+28 * -3.4128537e+22 = -3.5570482e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000001001000110011110110000;
		b = 32'b10011000000101100110111101110011;
		correct = 32'b01110000001001000110011110110000;
		#400 //2.0352357e+29 * -1.9443313e-24 = 2.0352357e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101110001010001010000101111;
		b = 32'b00010001111101110011101101100000;
		correct = 32'b00010001111101110011101101100001;
		#400 //1.8533205e-35 * 3.9006321e-28 = 3.9006324e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110100001110010100101001110;
		b = 32'b10010000100100101010110111000011;
		correct = 32'b00100110100001110010100101001110;
		#400 //9.378702e-16 * -5.785457e-29 = 9.378702e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010011100010010001111110110;
		b = 32'b10101100101011101110111110111111;
		correct = 32'b10111010011100010010001111110110;
		#400 //-0.0009198779 * -4.9719946e-12 = -0.0009198779
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000100000010111011001110110;
		b = 32'b11100011100001101101111101001110;
		correct = 32'b11100011100001101101111101010000;
		#400 //-1138766300000000.0 * -4.975909e+21 = -4.97591e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000010011100011010100010000;
		b = 32'b01010101111111110100001100111011;
		correct = 32'b01010101111111110100001100111011;
		#400 //211156.25 * 35083027000000.0 = 35083027000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001111011100100110111111100;
		b = 32'b10110001010010000111101110110011;
		correct = 32'b01001001111011100100110111111100;
		#400 //1952191.5 * -2.9174145e-09 = 1952191.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100010100110000010101101000;
		b = 32'b11010100011101000110100101101111;
		correct = 32'b11010100111000111011011101101100;
		#400 //-3625315200000.0 * -4198963600000.0 = -7824279000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001111101100011110111101111;
		b = 32'b00110011000110010100101001111110;
		correct = 32'b11001001111101100011110111101111;
		#400 //-2017213.9 * 3.569084e-08 = -2017213.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111000000000000100110000011;
		b = 32'b10101101011111011011011001010011;
		correct = 32'b11010111000000000000100110000011;
		#400 //-140778340000000.0 * -1.4421869e-11 = -140778340000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011011010000001100000111011;
		b = 32'b00100010100000100100001010000110;
		correct = 32'b11111011011010000001100000111011;
		#400 //-1.2051043e+36 * 3.5307005e-18 = -1.2051043e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001001100110011101111000100;
		b = 32'b11101110111111000001111001000100;
		correct = 32'b11101110111111000001111001000100;
		#400 //9.266153e-24 * -3.9013406e+28 = -3.9013406e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101000010011001010000110001;
		b = 32'b11101011011110110000110000110101;
		correct = 32'b11101011011110110000110000110101;
		#400 //-6.1960016e+17 * -3.0349803e+26 = -3.0349803e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100100001101001001010000101;
		b = 32'b10100100110000001110000001010000;
		correct = 32'b10111100100001101001001010000101;
		#400 //-0.016427288 * -8.364673e-17 = -0.016427288
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011111110100010010010111000;
		b = 32'b11011100111100011011001111001101;
		correct = 32'b11011100111100011011001111001101;
		#400 //-1.470211e-36 * -5.442653e+17 = -5.442653e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111111110011101000000000111;
		b = 32'b11010110101010011011000000111110;
		correct = 32'b11101111111110011101000000000111;
		#400 //-1.5462651e+29 * -93287210000000.0 = -1.5462651e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110001110101100001011000011;
		b = 32'b00001011100101001101010111010000;
		correct = 32'b01011110001110101100001011000011;
		#400 //3.3643833e+18 * 5.7329236e-32 = 3.3643833e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100111011011010100110000111;
		b = 32'b11010101011110110000101001100100;
		correct = 32'b01101100111011011010100110000111;
		#400 //2.2985279e+27 * -17251378000000.0 = 2.2985279e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011001001100111011000110110;
		b = 32'b00101111111011000100001110110000;
		correct = 32'b11111011001001100111011000110110;
		#400 //-8.643189e+35 * 4.2976245e-10 = -8.643189e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110101001000100011100110010;
		b = 32'b11010001101011110001011101101100;
		correct = 32'b11010001101011110001011101101100;
		#400 //2.654056e-25 * -94001530000.0 = -94001530000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101011011110001101011101110;
		b = 32'b01001100111100011010100100101101;
		correct = 32'b01001100111100011010100100101101;
		#400 //2.073907e-16 * 126699880.0 = 126699880.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110110100111101001101110000;
		b = 32'b11101101011010001010100110001101;
		correct = 32'b11101101011010001010100110001101;
		#400 //7.968006e-35 * -4.5003435e+27 = -4.5003435e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001101110100111111011001001;
		b = 32'b11111000000110100001000111011010;
		correct = 32'b11111000000110100001000111011010;
		#400 //1.263741e-18 * -1.2499622e+34 = -1.2499622e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011000011011010111110011011;
		b = 32'b11001100011010010000101100111000;
		correct = 32'b01110011000011011010111110011011;
		#400 //1.1225518e+31 * -61091040.0 = 1.1225518e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010111001101111111001100111;
		b = 32'b01111011111101011010000111111100;
		correct = 32'b01111011111101011010000111111100;
		#400 //6.2610984e-18 * 2.5507963e+36 = 2.5507963e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110110011110111000010001010;
		b = 32'b00010111010010000101011010001100;
		correct = 32'b11111110110011110111000010001010;
		#400 //-1.3786727e+38 * 6.4732723e-25 = -1.3786727e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111101100101001110010110111;
		b = 32'b00111001011000001001001110000010;
		correct = 32'b00111001011101101110011100011001;
		#400 //2.129223e-05 * 0.00021417256 = 0.00023546479
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101101000100000111101110010;
		b = 32'b01101011001111010100101110001000;
		correct = 32'b01101101101001111111100111001110;
		#400 //6.2694055e+27 * 2.2884367e+26 = 6.498249e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000011101111011110110110000;
		b = 32'b01001100101010101010000000110001;
		correct = 32'b01001100101010101010000000110001;
		#400 //4.885829e-29 * 89457030.0 = 89457030.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100100100110011110111001000;
		b = 32'b10101001110110101101100010001011;
		correct = 32'b10101001110110101101100010001011;
		#400 //-9.743614e-22 * -9.718709e-14 = -9.718709e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000011111011110000011101111;
		b = 32'b00110010101001010110000001010010;
		correct = 32'b01001000011111011110000011101111;
		#400 //259971.73 * 1.925233e-08 = 259971.73
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000101011010111101001001000;
		b = 32'b11100110010111000011010110110011;
		correct = 32'b11100110010111000011010110110011;
		#400 //6.842487e-29 * -2.599778e+23 = -2.599778e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100000101010111100101011011;
		b = 32'b00100101011101110111000010101001;
		correct = 32'b01011100000101010111100101011011;
		#400 //1.6829281e+17 * 2.1462006e-16 = 1.6829281e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111000000011110000110000010;
		b = 32'b10000001111101010000011000011010;
		correct = 32'b00111111000000011110000110000010;
		#400 //0.5073472 * -9.000754e-38 = 0.5073472
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101110000001010100000000010;
		b = 32'b11101010101011010100100001011101;
		correct = 32'b11101010101011010100100001011101;
		#400 //-1.811731e-35 * -1.0474295e+26 = -1.0474295e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110010010111010011010000000;
		b = 32'b00100001111111010010011111000110;
		correct = 32'b01010110010010111010011010000000;
		#400 //55978993000000.0 * 1.7154475e-18 = 55978993000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000000101101100011001111111;
		b = 32'b01010101011001000110000100001010;
		correct = 32'b01010101011001000110000100001010;
		#400 //-2.97352e-29 * 15694089000000.0 = 15694089000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011110100011000101001111101;
		b = 32'b11000001010101000111111011010101;
		correct = 32'b11000001010101000111111011010101;
		#400 //-9.757512e-08 * -13.280965 = -13.280965
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111000111101110001110011010;
		b = 32'b01010111000010101111011110010001;
		correct = 32'b01100111000111101110001110011010;
		#400 //7.503324e+23 * 152795900000000.0 = 7.503324e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001101101111001100000011000;
		b = 32'b00100100011101011110011110101001;
		correct = 32'b00101001101101111011011011010101;
		#400 //8.1532166e-14 * 5.332213e-17 = 8.158549e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100011101000101101101111101011;
		b = 32'b11110011110100000011001111111000;
		correct = 32'b11110011110100000011001111111000;
		#400 //-1.7657214e-17 * -3.2991083e+31 = -3.2991083e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111110101101100110110001111;
		b = 32'b11101110000111110110010110101011;
		correct = 32'b01111111110101101100110110001111;
		#400 //nan * -1.2332756e+28 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011110011111110001100010101;
		b = 32'b00011010101011111011011011100101;
		correct = 32'b00111011110011111110001100010101;
		#400 //0.006344209 * 7.2673786e-23 = 0.006344209
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011110111001010100101010010;
		b = 32'b01001111000010011000101101011000;
		correct = 32'b01001111000010011000101101011000;
		#400 //2.3924158e-17 * 2307610600.0 = 2307610600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000001000011100101100110011;
		b = 32'b11101101010100111101110101101010;
		correct = 32'b11101101010100111101110101101010;
		#400 //2.5280273 * -4.098063e+27 = -4.098063e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111000100001000001100101010111;
		b = 32'b01001111101001101101111001100001;
		correct = 32'b01111000100001000001100101010111;
		#400 //2.1434286e+34 * 5599183400.0 = 2.1434286e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111000011100001011010100011;
		b = 32'b10000000011101110111001001010101;
		correct = 32'b01111111000011100001011010100011;
		#400 //1.8886791e+38 * -1.0969439e-38 = 1.8886791e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100011101010000000010100111;
		b = 32'b01011011111011011111101010101011;
		correct = 32'b01011011111011011111101010101011;
		#400 //980.0102 * 1.3397036e+17 = 1.3397036e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101010000100110000110001111;
		b = 32'b10011100000111100000100110010100;
		correct = 32'b00011101000110101101111100101010;
		#400 //2.5726123e-21 * -5.2290194e-22 = 2.0497103e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100100100100111000110000111;
		b = 32'b00110011010010010011101101000110;
		correct = 32'b01001100100100100111000110000111;
		#400 //76778550.0 * 4.685287e-08 = 76778550.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110011011100111100100110111;
		b = 32'b00110101011011000111000111010101;
		correct = 32'b01111110011011100111100100110111;
		#400 //7.924641e+37 * 8.80825e-07 = 7.924641e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101110110100100111110011011;
		b = 32'b11001000011010011100011100000010;
		correct = 32'b11001000011010011100011100000010;
		#400 //-5.778643e-21 * -239388.03 = -239388.03
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001101100101101001011111010;
		b = 32'b11000011000000000001110001100101;
		correct = 32'b11000011000000000001110001100101;
		#400 //-4.3050343e-33 * -128.11092 = -128.11092
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000000011110101101001001001;
		b = 32'b11001011000000010110111101000110;
		correct = 32'b01010000000011110011100111101101;
		#400 //9620235000.0 * -8482630.0 = 9611752000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111101011010111101000100010;
		b = 32'b10100110011000101001010010111111;
		correct = 32'b10110111101011010111101000100010;
		#400 //-2.068008e-05 * -7.861109e-16 = -2.068008e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000011100010100001110000100;
		b = 32'b10000010100111000001110110010000;
		correct = 32'b11010000011100010100001110000100;
		#400 //-16190935000.0 * -2.2939108e-37 = -16190935000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111110101111000010010110010;
		b = 32'b11100011110111110000110001010100;
		correct = 32'b11111111110101111000010010110010;
		#400 //nan * -8.2290245e+21 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011010111000101111010001110;
		b = 32'b00001010101000000110010000011001;
		correct = 32'b01101011010111000101111010001110;
		#400 //2.664102e+26 * 1.5445092e-32 = 2.664102e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111001001111000111000101110;
		b = 32'b00101001110100000111110110011010;
		correct = 32'b00101001110100000111110110011010;
		#400 //1.2605466e-34 * 9.258844e-14 = 9.258844e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001100110111100011000111110;
		b = 32'b01110100110011001100101100111010;
		correct = 32'b11111001100110111001001100001011;
		#400 //-1.0110336e+35 * 1.2980353e+32 = -1.0097355e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101101001000000011011001111;
		b = 32'b01110101000101000110111101111111;
		correct = 32'b01110101000101000110111101111111;
		#400 //1.5424987e-35 * 1.881644e+32 = 1.881644e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011111101001101010010010100;
		b = 32'b00010110000101000100111001010101;
		correct = 32'b11011011111101001101010010010100;
		#400 //-1.3782725e+17 * 1.1980062e-25 = -1.3782725e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010011110111111110111000110;
		b = 32'b11010110001100110011101001001111;
		correct = 32'b11010110001100110011101001001111;
		#400 //-2.2381324e-13 * -49265754000000.0 = -49265754000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001001111000011101110000101;
		b = 32'b11101011011010110001011001011001;
		correct = 32'b11101011011010110001011001011001;
		#400 //2.2657663e-33 * -2.842031e+26 = -2.842031e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011011101110000001101001010;
		b = 32'b01111011110111010100011010001110;
		correct = 32'b01111011010000111000100111010010;
		#400 //-1.282564e+36 * 2.2978572e+36 = 1.0152932e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000111011001111001010111101;
		b = 32'b10111000100000100100100100011001;
		correct = 32'b11010000111011001111001010111101;
		#400 //-31802649000.0 * -6.2124986e-05 = -31802649000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010101000000111111111001111110;
		b = 32'b10100000011111000100101111000001;
		correct = 32'b10100000011111000100101111000011;
		#400 //-2.6655998e-26 * -2.1370295e-19 = -2.1370298e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111100011000010011011110111;
		b = 32'b10100100011001010100001100100110;
		correct = 32'b10100100011001010100001100100110;
		#400 //1.3820075e-29 * -4.9713336e-17 = -4.9713336e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101010110100001011000000110;
		b = 32'b11001111011010100110000010100011;
		correct = 32'b11001111010111001011111101000011;
		#400 //228679780.0 * -3932201700.0 = -3703522000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001110001010011110000100110;
		b = 32'b11101111011110111001000100000111;
		correct = 32'b11101111011110111001000100000111;
		#400 //-4.748259e-33 * -7.7856065e+28 = -7.7856065e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101000111000101101111000111;
		b = 32'b11010100100100011101010110100010;
		correct = 32'b11111101000111000101101111000111;
		#400 //-1.2989756e+37 * -5010835400000.0 = -1.2989756e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010010000010001101110110011001;
		b = 32'b10001110100000001111100000011101;
		correct = 32'b00010010000001111101101110101001;
		#400 //4.3187173e-28 * -3.179336e-30 = 4.286924e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011101011001101011101100000;
		b = 32'b00100000010001110100100110001110;
		correct = 32'b00100000010001111001111111111010;
		#400 //2.8594196e-22 * 1.6880293e-19 = 1.6908887e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100000111110000110111010010;
		b = 32'b11011001110001011111010111001001;
		correct = 32'b11011001110001011111010111001001;
		#400 //0.009707885 * -6965102000000000.0 = -6965102000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110001111000010110001001001;
		b = 32'b11011111111111011101101110001111;
		correct = 32'b11011111111111011101101110001111;
		#400 //-9.961795e-21 * -3.6584743e+19 = -3.6584743e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010011101111010000001011011;
		b = 32'b00010001100001001010010100101001;
		correct = 32'b01100010011101111010000001011011;
		#400 //1.14197515e+21 * 2.0927716e-28 = 1.14197515e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001110110001110110001101110111;
		b = 32'b11101100110110101001000101010111;
		correct = 32'b11101100110110101001000101010111;
		#400 //1672592300.0 * -2.1138574e+27 = -2.1138574e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100111111110111111100111000;
		b = 32'b01100010101001101000111001110111;
		correct = 32'b11111100111111110111111100111000;
		#400 //-1.0612928e+37 * 1.5362126e+21 = -1.0612928e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111101101100010010001000101;
		b = 32'b11000110000110101001011111111011;
		correct = 32'b11010111101101100010010001000101;
		#400 //-400533800000000.0 * -9893.995 = -400533800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011101011101110001001101100;
		b = 32'b01101111101011101011011101111001;
		correct = 32'b01101111101011101011011101111001;
		#400 //-1502246100000.0 * 1.0814439e+29 = 1.0814439e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110101100110111001111010011;
		b = 32'b00000110110110100001010111000101;
		correct = 32'b00100110101100110111001111010011;
		#400 //1.2452014e-15 * 8.2034473e-35 = 1.2452014e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101111011010000111010011001;
		b = 32'b10001010011111100110010110000100;
		correct = 32'b01001101111011010000111010011001;
		#400 //497144600.0 * -1.2248748e-32 = 497144600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101000010100001001001000110;
		b = 32'b00100101110001110000111010110000;
		correct = 32'b01100101000010100001001001000110;
		#400 //4.075148e+22 * 3.453095e-16 = 4.075148e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011001101100011010100000011;
		b = 32'b10011111001100010111110011010010;
		correct = 32'b00110011001101100011010100000011;
		#400 //4.242339e-08 * -3.7584457e-20 = 4.242339e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001010111101010100000110101;
		b = 32'b00111100000101110001010000000100;
		correct = 32'b00111100000101110001010000000100;
		#400 //-4.0895643e-38 * 0.009221081 = 0.009221081
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001110010000011011110110011;
		b = 32'b00001101001011010001111001001101;
		correct = 32'b10110001110010000011011110110011;
		#400 //-5.8270984e-09 * 5.3346214e-31 = -5.8270984e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011000011100010011110100011;
		b = 32'b10010100000110001101010101100011;
		correct = 32'b01001011000011100010011110100011;
		#400 //9316259.0 * -7.716122e-27 = 9316259.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100110101000001101100010001;
		b = 32'b11010101101110011110001010001110;
		correct = 32'b11010101101110011110001010001110;
		#400 //-1.403598e-21 * -25547837000000.0 = -25547837000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000000001011111110100110001;
		b = 32'b11011111001011011001110000011010;
		correct = 32'b11011111001011011001110000011010;
		#400 //-2.0935786 * -1.2509902e+19 = -1.2509902e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001010001011100010100001000;
		b = 32'b01110000101101010000111101011111;
		correct = 32'b01110000101101010000111101011111;
		#400 //12.360603 * 4.4828295e+29 = 4.4828295e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100110001100111000101111010;
		b = 32'b01111000010111001001010000111011;
		correct = 32'b01111000010111001001010000111101;
		#400 //1.9192255e+27 * 1.7895497e+34 = 1.7895499e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000000110010011111010000001;
		b = 32'b11000110100010001111111000100101;
		correct = 32'b11000110100010001111111000100101;
		#400 //-1.2980285e-19 * -17535.072 = -17535.072
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000001111011101101111010110;
		b = 32'b11001000000011001010111011111100;
		correct = 32'b11001000000011001010111011111100;
		#400 //5.7133535e-34 * -144059.94 = -144059.94
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011111100100100000000101010;
		b = 32'b11000111000011001110100001100010;
		correct = 32'b11111011111100100100000000101010;
		#400 //-2.5156745e+36 * -36072.383 = -2.5156745e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110010110001001010011011010;
		b = 32'b01010101111110010011010111001110;
		correct = 32'b01100110010110001001010011011010;
		#400 //2.5569425e+23 * 34251186000000.0 = 2.5569425e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101100010001000011100010110;
		b = 32'b10011011101111001110101010000111;
		correct = 32'b01011101100010001000011100010110;
		#400 //1.229732e+18 * -3.125355e-22 = 1.229732e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101111000111010111100010100000;
		b = 32'b10010010010110011101001110100111;
		correct = 32'b00101111000111010111100010100000;
		#400 //1.4321921e-10 * -6.873401e-28 = 1.4321921e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010100100001001111000110000;
		b = 32'b11101010101010000101101101001001;
		correct = 32'b11101010101010000101101101001001;
		#400 //5.981257e-23 * -1.0176531e+26 = -1.0176531e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000000100101110000110010000;
		b = 32'b11011111001001110011000001001101;
		correct = 32'b11011111001001110011000001001101;
		#400 //5.3435034e-10 * -1.2047214e+19 = -1.2047214e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110011011011001011000101000;
		b = 32'b10101010000111111000011010101101;
		correct = 32'b10101010000111111000011010101101;
		#400 //-1.9192088e-25 * -1.4168762e-13 = -1.4168762e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101110000011011000011110100;
		b = 32'b00011110001010001001111110110101;
		correct = 32'b11001101110000011011000011110100;
		#400 //-406199940.0 * 8.9268726e-21 = -406199940.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100100111101000101010110100;
		b = 32'b01100011100100010111110000000011;
		correct = 32'b11100100011101000101011101100110;
		#400 //-2.3396641e+22 * 5.367428e+21 = -1.8029213e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111110110111100110001000010;
		b = 32'b10111101110110101101010110110110;
		correct = 32'b11011111110110111100110001000010;
		#400 //-3.1676213e+19 * -0.106852934 = -3.1676213e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011011000000111110011000001;
		b = 32'b01110000111000101111110101010010;
		correct = 32'b01110000111000101111110101010010;
		#400 //224.48732 * 5.6199886e+29 = 5.6199886e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001111101000001110000100000;
		b = 32'b10101111100100011000111110001101;
		correct = 32'b10101111100100011000111110001101;
		#400 //2.5240368e-23 * -2.6477345e-10 = -2.6477345e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111100010100010101100001001;
		b = 32'b11001111100001011110111000100011;
		correct = 32'b01011111100010100010101100001001;
		#400 //1.9912123e+19 * -4493952500.0 = 1.9912123e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110001110100110011101000000;
		b = 32'b01000111010110100110011111001111;
		correct = 32'b11010110001110100110011101000000;
		#400 //-51238155000000.0 * 55911.81 = -51238155000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000010110011110101110100101;
		b = 32'b11101110110011100111100101111101;
		correct = 32'b11101110110011100111100101111101;
		#400 //-223150.58 * -3.195039e+28 = -3.195039e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010000001111001010110111111;
		b = 32'b01010000010001110111101011101110;
		correct = 32'b01010000010001110111101011101110;
		#400 //-7.8920825e-09 * 13386889000.0 = 13386889000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011010011101100011110101110;
		b = 32'b11001011101010001011100110011001;
		correct = 32'b11111011010011101100011110101110;
		#400 //-1.0736631e+36 * -22115122.0 = -1.0736631e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100001000000001011111001001;
		b = 32'b11011000101001010011000100100111;
		correct = 32'b11011000101001010011000100100111;
		#400 //3.4714616e-17 * -1453044200000000.0 = -1453044200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010100000011101010010111000;
		b = 32'b10110010100110001000100111000001;
		correct = 32'b10110001001101011010100001001000;
		#400 //1.511431e-08 * -1.7757772e-08 = -2.6434623e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110101000101111101011001011;
		b = 32'b00011001110101100111001100110101;
		correct = 32'b11110110101000101111101011001011;
		#400 //-1.6528101e+33 * 2.2173613e-23 = -1.6528101e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001011001000010111000001100;
		b = 32'b01101001001010011110001110001000;
		correct = 32'b11101000011010010010101000010000;
		#400 //-1.7240784e+25 * 1.2836434e+25 = -4.4043492e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111000011111101110110010111;
		b = 32'b10110010100100111100000011101010;
		correct = 32'b10110010100100111100000011101010;
		#400 //-7.093121e-30 * -1.720078e-08 = -1.720078e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000000001000010100111001000;
		b = 32'b01101011111101110001100001101010;
		correct = 32'b01101011111101110001100001101010;
		#400 //8869323000.0 * 5.9743994e+26 = 5.9743994e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010111100010110110110010111;
		b = 32'b00110111001001111110101101010111;
		correct = 32'b00110111001001111110101101010111;
		#400 //6.5439214e-18 * 1.000877e-05 = 1.000877e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101001101001011100001101101;
		b = 32'b01101100100000000010010101111010;
		correct = 32'b01101101011101001100101100101010;
		#400 //3.4956412e+27 * 1.2393559e+27 = 4.734997e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011111100111101100110001000;
		b = 32'b00100010110110011111101010010100;
		correct = 32'b01100011111100111101100110001000;
		#400 //8.996467e+21 * 5.9083278e-18 = 8.996467e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111010001110101001101000001;
		b = 32'b10111110011101101010001111111111;
		correct = 32'b11101111010001110101001101000001;
		#400 //-6.1688165e+28 * -0.24085997 = -6.1688165e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101010011010001001010110111;
		b = 32'b00011000001110011001110101011111;
		correct = 32'b11101101010011010001001010110111;
		#400 //-3.9666907e+27 * 2.3990142e-24 = -3.9666907e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000001100010001000011100010;
		b = 32'b01001100011011000111100100001100;
		correct = 32'b01100000001100010001000011100010;
		#400 //5.1035785e+19 * 61989936.0 = 5.1035785e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011001000110110001100000001;
		b = 32'b00000110110000001011101011000110;
		correct = 32'b00111011001000110110001100000001;
		#400 //0.0024930837 * 7.249681e-35 = 0.0024930837
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101111000111111011101000001;
		b = 32'b10100100101100100110001101100010;
		correct = 32'b11001101111000111111011101000001;
		#400 //-478079000.0 * -7.7363556e-17 = -478079000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000101010111010000001001000;
		b = 32'b10010010010010110101110111101100;
		correct = 32'b11101000101010111010000001001000;
		#400 //-6.4838507e+24 * -6.4171273e-28 = -6.4838507e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000101010011100011001100100;
		b = 32'b01110000001110010100000101011010;
		correct = 32'b11110000000110100100101101101110;
		#400 //-4.2034245e+29 * 2.2933493e+29 = -1.9100752e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001110011000010100100011100;
		b = 32'b00100000000000000110111001100000;
		correct = 32'b00100000000000000110111001100000;
		#400 //-7.4996754e-38 * 1.0878542e-19 = 1.0878542e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110110011101011110011010100;
		b = 32'b10011010101010101001000011110001;
		correct = 32'b00100110110011101011110011010011;
		#400 //1.4345303e-15 * -7.054452e-23 = 1.4345302e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001111010010000011110011010;
		b = 32'b01110000010110111100001011000110;
		correct = 32'b01111001111010010000011110110101;
		#400 //1.5124492e+35 * 2.7205074e+29 = 1.5124519e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101111010000011111011101100;
		b = 32'b00101001001111001111101100001001;
		correct = 32'b00101001001111001111101100001011;
		#400 //6.147495e-21 * 4.1962124e-14 = 4.196213e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001110011110010001011000001110;
		b = 32'b11001110000110011101000010110001;
		correct = 32'b01001101101111101000101010111010;
		#400 //1044743040.0 * -645147700.0 = 399595330.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000000100100101001100100100;
		b = 32'b11011000000010000101011111101001;
		correct = 32'b11011000000010000101011111101001;
		#400 //4.403301e-34 * -599644600000000.0 = -599644600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010100110010001010010010111;
		b = 32'b10111101111110000010010111111000;
		correct = 32'b10111101111110000010010111111000;
		#400 //6.331258e-23 * -0.12116617 = -0.12116617
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001110000111010011001011010010;
		b = 32'b00110100110010100101101010110111;
		correct = 32'b00110100110010100101101010110111;
		#400 //1.9376213e-30 * 3.7691436e-07 = 3.7691436e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111001101000010101010101111;
		b = 32'b00110100101110111110111100110001;
		correct = 32'b00110100101110111110111100110001;
		#400 //1.3554239e-34 * 3.50055e-07 = 3.50055e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000000111111001010100010011;
		b = 32'b00100011000000001100000111101011;
		correct = 32'b00100011000000110100000000111111;
		#400 //1.3517148e-19 * 6.979958e-18 = 7.115129e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010000011110101111000100000;
		b = 32'b00000010011100110100101010110100;
		correct = 32'b00001010000011110101111100010011;
		#400 //6.9029025e-33 * 1.7874259e-37 = 6.903081e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110101111011011000111001010;
		b = 32'b00101011000110010011001011011111;
		correct = 32'b11001110101111011011000111001010;
		#400 //-1591272700.0 * 5.4427117e-13 = -1591272700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101010101100100010011001110;
		b = 32'b10000111100001111110010110001011;
		correct = 32'b11001101010101100100010011001110;
		#400 //-224677090.0 * -2.0447456e-34 = -224677090.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111010100101111010111011111;
		b = 32'b11011000010001010111111000010000;
		correct = 32'b11011000010001010111111000010000;
		#400 //54005.87 * -868580900000000.0 = -868580900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101111110101011000110101001101;
		b = 32'b11111100011001000001101000011101;
		correct = 32'b11111100011001000001101000011101;
		#400 //3.8844875e-10 * -4.7374933e+36 = -4.7374933e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000111011100100100100111110;
		b = 32'b01010110010101001011010110101011;
		correct = 32'b01100000111011100100100101000101;
		#400 //1.3736259e+20 * 58469180000000.0 = 1.3736265e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010011000000100100000100001;
		b = 32'b00010100010001011111111000101010;
		correct = 32'b10101010011000000100100000100001;
		#400 //-1.9920221e-13 * 9.996083e-27 = -1.9920221e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010010000110010000001011100;
		b = 32'b10001100000101000111101010000010;
		correct = 32'b11001010010000110010000001011100;
		#400 //-3196951.0 * -1.1438371e-31 = -3196951.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000000010000000001110111001;
		b = 32'b10100111010110101100111111111001;
		correct = 32'b10100111010110101100111111111001;
		#400 //-7.3602e-40 * -3.036632e-15 = -3.036632e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001000000110111101110101001;
		b = 32'b00011011011010110111001010110111;
		correct = 32'b11001001000000110111101110101001;
		#400 //-538554.56 * 1.9475811e-22 = -538554.56
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100101111110001010011110101;
		b = 32'b01001101010010110110000101110011;
		correct = 32'b01001101010010110110000101110011;
		#400 //8.286855e-17 * 213260080.0 = 213260080.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010110100000001010100011000;
		b = 32'b01001011010010000101110011011100;
		correct = 32'b01001011010010000101110011011100;
		#400 //-2.422398e-08 * 13130972.0 = 13130972.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110010101001101101110111101;
		b = 32'b11010111001110000000011010110001;
		correct = 32'b11100110010101001101101110111101;
		#400 //-2.5129879e+23 * -202338880000000.0 = -2.5129879e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100111101000011011001010101;
		b = 32'b00100100010001000101101000110100;
		correct = 32'b00110100111101000011011001010101;
		#400 //4.5488073e-07 * 4.257713e-17 = 4.5488073e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000011100000101001100111110;
		b = 32'b00001001110100110010001101101000;
		correct = 32'b11000000011100000101001100111110;
		#400 //-3.7550807 * 5.0829698e-33 = -3.7550807
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010110000011110100110100001;
		b = 32'b01111100101101111111100111001011;
		correct = 32'b01111100101101111111100111001011;
		#400 //-8.020038e-23 * 7.642054e+36 = 7.642054e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010111101100110000101010010;
		b = 32'b00110011000110000110010011101011;
		correct = 32'b01001010111101100110000101010010;
		#400 //8073385.0 * 3.5482042e-08 = 8073385.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000010000100100110100011010;
		b = 32'b01100111110001110100010011011011;
		correct = 32'b01100111110001110100010011011011;
		#400 //-198964.4 * 1.8820422e+24 = 1.8820422e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100001101010100011000110011;
		b = 32'b11100000101001100100101010111101;
		correct = 32'b11100000101001100100101010111101;
		#400 //3.930758e-17 * -9.586078e+19 = -9.586078e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010101111101110001001101000;
		b = 32'b01110111011100011110011010010011;
		correct = 32'b01110111011100011110011010010011;
		#400 //-6254900.0 * 4.9063287e+33 = 4.9063287e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111100111100101101000011001;
		b = 32'b01100111101011101001010101100100;
		correct = 32'b01100111101011101001010101100100;
		#400 //81076.195 * 1.6488951e+24 = 1.6488951e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100100110101011101110100001001;
		b = 32'b11010100100011000001100011000001;
		correct = 32'b11010100100011000001100011000001;
		#400 //-9.274847e-17 * -4813686000000.0 = -4813686000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011010000101010101010101000;
		b = 32'b10000010001000010000100100100011;
		correct = 32'b00100011010000101010101010101000;
		#400 //1.0552899e-17 * -1.1831034e-37 = 1.0552899e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000001010011110111110100000;
		b = 32'b11010011001101110011011110110101;
		correct = 32'b11010011001110011101111101110100;
		#400 //-11404214000.0 * -786913600000.0 = -798317900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000011000111011111010110100;
		b = 32'b11011001100000010011100101100101;
		correct = 32'b11011001100000010011100101100101;
		#400 //-5.4298624e-05 * -4546672000000000.0 = -4546672000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010011010001111010111111001;
		b = 32'b10100101111010111110111000110011;
		correct = 32'b01011010011010001111010111111001;
		#400 //1.6393161e+16 * -4.0927412e-16 = 1.6393161e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101110011111001110101010000;
		b = 32'b10001000000110011000110001111110;
		correct = 32'b11100101110011111001110101010000;
		#400 //-1.2255397e+23 * -4.620691e-34 = -1.2255397e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011100010111000000000010000;
		b = 32'b11000111011100001011110100011110;
		correct = 32'b11000111011100001011110100011110;
		#400 //2.307838e-22 * -61629.117 = -61629.117
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010011110001010110001011101;
		b = 32'b00001010111011011110001111110001;
		correct = 32'b11110010011110001010110001011101;
		#400 //-4.925482e+30 * 2.2908012e-32 = -4.925482e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101010011110110101100000001;
		b = 32'b01100011111111101111010001111100;
		correct = 32'b01100011111111101111010001111100;
		#400 //-7.726922e-07 * 9.40618e+21 = 9.40618e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111001101010100010011101000;
		b = 32'b01000100000111000110101111000111;
		correct = 32'b01000100000111000011111001110110;
		#400 //-0.7080827 * 625.684 = 624.97595
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101101001001111100001011110;
		b = 32'b01010100100101001110100011111101;
		correct = 32'b11010101011111110111110000111110;
		#400 //-22673330000000.0 * 5116512400000.0 = -17556818000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001010010001101101101010010;
		b = 32'b10000111111101101001010101010010;
		correct = 32'b00001001001010100000100010101000;
		#400 //2.4177248e-33 * -3.7101729e-34 = 2.0467076e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000100111111000100111011111;
		b = 32'b01110111011011000010101111011110;
		correct = 32'b01110111011011000010101111011110;
		#400 //4.98558 * 4.7901242e+33 = 4.7901242e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011101000001100100010101111;
		b = 32'b10000000111010111101010100011110;
		correct = 32'b10101011101000001100100010101111;
		#400 //-1.1424385e-12 * -2.1657794e-38 = -1.1424385e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111100100001110111111001100;
		b = 32'b11100011000111000010101010111100;
		correct = 32'b11100011000111000010101010111100;
		#400 //-4863269000.0 * -2.8807714e+21 = -2.8807714e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111000001010010010100010010100;
		b = 32'b01101011101101111010001100110000;
		correct = 32'b01111000001010010010100010010100;
		#400 //1.3723769e+34 * 4.440081e+26 = 1.3723769e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010010101110011010000010001;
		b = 32'b01100000111000011000100111101100;
		correct = 32'b01110010010101110011010000010001;
		#400 //4.2625422e+30 * 1.3001424e+20 = 4.2625422e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110110001000010001110100101;
		b = 32'b11001011011111000010000111011101;
		correct = 32'b11001011011111000010000111011101;
		#400 //-1.3609894e-15 * -16523741.0 = -16523741.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111111101111010110001111001;
		b = 32'b11100011110010110011100101111001;
		correct = 32'b11100011110010110011100101111001;
		#400 //1.6005539e-24 * -7.497661e+21 = -7.497661e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010110000011001000001100001;
		b = 32'b11001101000010100100100010100100;
		correct = 32'b11110010110000011001000001100001;
		#400 //-7.667859e+30 * -145001020.0 = -7.667859e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111010011111011000001100010000;
		b = 32'b11100100100010000011011100110011;
		correct = 32'b11100100100010000011011100110011;
		#400 //0.0009670714 * -2.0101878e+22 = -2.0101878e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011010110111110100000011001;
		b = 32'b10001101001110111011010100111001;
		correct = 32'b00110011010110111110100000011001;
		#400 //5.1201003e-08 * -5.7841963e-31 = 5.1201003e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100000101010111110011011100;
		b = 32'b11100001111111100011010110111111;
		correct = 32'b01100100000011011000101100101110;
		#400 //1.1030248e+22 * -5.8616823e+20 = 1.044408e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111011100100111111111101110;
		b = 32'b10011100111000010110110001000011;
		correct = 32'b01000111011100100111111111101110;
		#400 //62079.93 * -1.4917236e-21 = 62079.93
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111100100111010111111000111;
		b = 32'b00101000110101001011011110111101;
		correct = 32'b00101000111110011010001110101111;
		#400 //4.0991274e-15 * 2.3616412e-14 = 2.771554e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110101100010011000011101001;
		b = 32'b01001001111101010011000101101101;
		correct = 32'b01001001111101010011000101101101;
		#400 //-1.2295099e-15 * 2008621.6 = 2008621.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000111110101110111010000001;
		b = 32'b00101101010110101100001110100100;
		correct = 32'b11011000111110101110111010000001;
		#400 //-2207218200000000.0 * 1.2435306e-11 = -2207218200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001000001111101000100000001100;
		b = 32'b10001001100001001011000000101111;
		correct = 32'b10001001100111001000000100110000;
		#400 //-5.7335968e-34 * -3.1943526e-33 = -3.767712e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011111010011110001110100110;
		b = 32'b11111011010011110000100010000111;
		correct = 32'b11111011010011110000100010000111;
		#400 //-30656332.0 * -1.0749784e+36 = -1.0749784e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111010100010101100010001000;
		b = 32'b11010110100010011001011011110000;
		correct = 32'b11010110100010011001010101001101;
		#400 //3512240000.0 * -75640680000000.0 = -75637170000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011100010100001010010011001110;
		b = 32'b01010001001101100011110100010010;
		correct = 32'b01010001001101100011110100010010;
		#400 //6.903443e-22 * 48919290000.0 = 48919290000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101100101001011110110101100110;
		b = 32'b01001010010010011100100100110001;
		correct = 32'b01001010010010011100100100110001;
		#400 //4.7159386e-12 * 3306060.2 = 3306060.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001101000101111111000001010;
		b = 32'b01100100000111010010000111110110;
		correct = 32'b01100100000111010010000111110110;
		#400 //20.374043 * 1.1594344e+22 = 1.1594344e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010110110010001010111001000;
		b = 32'b00011001000111011100011101001001;
		correct = 32'b11000010110110010001010111001000;
		#400 //-108.54254 * 8.156955e-24 = -108.54254
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110010010001001011000011110;
		b = 32'b00011101101000010000010110001010;
		correct = 32'b01010110010010001001011000011110;
		#400 //55136770000000.0 * 4.2622072e-21 = 55136770000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111000010111100011101000000;
		b = 32'b11110001110001001100101000010011;
		correct = 32'b11110001110001001100101000010011;
		#400 //-2345091000.0 * -1.9489073e+30 = -1.9489073e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010111010001001101000100001;
		b = 32'b00011001100111011010010010100101;
		correct = 32'b00011001100111011010010010100101;
		#400 //3.4177802e-37 * 1.6299919e-23 = 1.6299919e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111010111001111110100011111;
		b = 32'b10011001110110111100011110111111;
		correct = 32'b10011001110110111100011111000110;
		#400 //-1.0895587e-29 * -2.2724746e-23 = -2.2724757e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011110010000101101001011110;
		b = 32'b00100010101111111101001000011101;
		correct = 32'b00100010101111111100111011111100;
		#400 //-3.3145623e-22 * 5.199312e-18 = 5.1989807e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101101011110010111000111110;
		b = 32'b11110001010100011111010100101110;
		correct = 32'b11110001010100011111010100101110;
		#400 //4.6369928e-21 * -1.0396603e+30 = -1.0396603e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100101010100111001001001101;
		b = 32'b00101001110101011101111100111011;
		correct = 32'b00110100101010100111001001010000;
		#400 //3.1748132e-07 * 9.4978245e-14 = 3.174814e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000101001011000011111101001;
		b = 32'b11010001111101000111011110101110;
		correct = 32'b11010001111101000111011110101110;
		#400 //6.529043e-29 * -131247490000.0 = -131247490000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100000101100010100100010010;
		b = 32'b00100001110100100110101110001111;
		correct = 32'b00100001110100100110101110001111;
		#400 //-7.581164e-27 * 1.4258624e-18 = 1.4258624e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110010010111010101100100100;
		b = 32'b10011111010101000101000110010101;
		correct = 32'b10100110010010111010111001110101;
		#400 //-7.066171e-16 * -4.496023e-20 = -7.0666206e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001010111100111001010100110;
		b = 32'b00001110100011010010110110101100;
		correct = 32'b01010001010111100111001010100110;
		#400 //59712890000.0 * 3.4803164e-30 = 59712890000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001011011001011010100101001;
		b = 32'b01101111001011010010000100011000;
		correct = 32'b01101111001011010010000100011000;
		#400 //3.4445498e-09 * 5.3580915e+28 = 5.3580915e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000011110000110110001011100;
		b = 32'b10010101000011111000011001111101;
		correct = 32'b10111000011110000110110001011100;
		#400 //-5.9228725e-05 * -2.8984713e-26 = -5.9228725e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011011111000001111011011001;
		b = 32'b10100111111111110111110110010111;
		correct = 32'b10100111111111110111110110010111;
		#400 //2.0854919e-22 * -7.0912883e-15 = -7.0912883e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011010000011000000100100011;
		b = 32'b10110010100101111010100111111011;
		correct = 32'b01011011010000011000000100100011;
		#400 //5.4466658e+16 * -1.7656012e-08 = 5.4466658e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111111001001010001100110000;
		b = 32'b00111010011101110110011110011001;
		correct = 32'b00111010011101110110011110011001;
		#400 //1.4775349e-24 * 0.00094377395 = 0.00094377395
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101100110101001011011010011;
		b = 32'b01100111000010100001000100111100;
		correct = 32'b01110101100110101001011011010011;
		#400 //3.9193008e+32 * 6.520045e+23 = 3.9193008e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000110110100111100010010000;
		b = 32'b10001110111011110010001100001111;
		correct = 32'b11110000110110100111100010010000;
		#400 //-5.4090787e+29 * -5.895181e-30 = -5.4090787e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111000010010110010001111101;
		b = 32'b10101000110001100010111110101011;
		correct = 32'b11010111000010010110010001111101;
		#400 //-151064690000000.0 * -2.2003089e-14 = -151064690000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000110000000111010111011001101;
		b = 32'b01001100110111010101100011100111;
		correct = 32'b01001100110111010101100011100111;
		#400 //-2.4766785e-35 * 116049720.0 = 116049720.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101100001101110011011100011;
		b = 32'b00110111110100110100011110010111;
		correct = 32'b01001101100001101110011011100011;
		#400 //282909800.0 * 2.5186497e-05 = 282909800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111100010110111111000100100;
		b = 32'b00011111110101000100101101100100;
		correct = 32'b01100111100010110111111000100100;
		#400 //1.3174716e+24 * 8.9910216e-20 = 1.3174716e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110001001111101011011100011;
		b = 32'b11111001111011111011011001011111;
		correct = 32'b11111001111011111011011001011111;
		#400 //-703969500.0 * -1.5558223e+35 = -1.5558223e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001010110000000000111010011;
		b = 32'b00001011001011100100011000101100;
		correct = 32'b01000001010110000000000111010011;
		#400 //13.500445 * 3.3563972e-32 = 13.500445
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011111101010010011000111110;
		b = 32'b10111110110111000010100100110111;
		correct = 32'b01101011111101010010011000111110;
		#400 //5.9273484e+26 * -0.43000194 = 5.9273484e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111110100111010010111110100;
		b = 32'b11100100010000010110001110100101;
		correct = 32'b11100100010000010110001110100101;
		#400 //1.3677448e-24 * -1.4269607e+22 = -1.4269607e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000001101011000111111101110;
		b = 32'b00110101001000101100000011001011;
		correct = 32'b10111000001100110000010011101011;
		#400 //-4.3287808e-05 * 6.0630254e-07 = -4.2681506e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011000000010011111111111111;
		b = 32'b00110101100010110001001100100001;
		correct = 32'b00110101100010110001001100100001;
		#400 //1.6313642e-27 * 1.0361874e-06 = 1.0361874e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101000010100001001000100000;
		b = 32'b10101011111100010011101011001100;
		correct = 32'b10111101000010100001001000100000;
		#400 //-0.03370869 * -1.7140399e-12 = -0.03370869
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001010001010111010011101111;
		b = 32'b11101101011010110110101111111101;
		correct = 32'b11101101011010110110101111111101;
		#400 //6.6900957e-19 * -4.5537204e+27 = -4.5537204e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111010001100011101001101001;
		b = 32'b01100010010000100000010000010010;
		correct = 32'b01100010010000100000010000010010;
		#400 //1.1815319e-05 * 8.947404e+20 = 8.947404e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100010010001010101110110000001;
		b = 32'b00001000100001101100111100101001;
		correct = 32'b11100010010001010101110110000001;
		#400 //-9.1018656e+20 * 8.113535e-34 = -9.1018656e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010110000001111111001111101;
		b = 32'b11001100011101001011111110010101;
		correct = 32'b01011010110000001111111001111101;
		#400 //2.7161504e+16 * -64159316.0 = 2.7161504e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010111100100010111101000111;
		b = 32'b10000001111010111110100111010000;
		correct = 32'b10001010111100100010111110000010;
		#400 //-2.3321536e-32 * -8.666087e-38 = -2.3321623e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110001110001101001010011100;
		b = 32'b10101111011110000111010010011101;
		correct = 32'b10111110001110001101001010011100;
		#400 //-0.18049091 * -2.2596898e-10 = -0.18049091
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111010001001010000100100110;
		b = 32'b11010100101011001110001010011000;
		correct = 32'b11010100101011001110001010011000;
		#400 //-0.76808393 * -5940288000000.0 = -5940288000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000110000111011111100101101;
		b = 32'b00110110001101110000111110010000;
		correct = 32'b00110110001101110000111110010000;
		#400 //-3.3160794e-19 * 2.7278184e-06 = 2.7278184e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110010001010111100101111001;
		b = 32'b00000011100000011011110000010010;
		correct = 32'b10110110010001010111100101111001;
		#400 //-2.9425994e-06 * 7.625117e-37 = -2.9425994e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101010010011000011110010000011;
		b = 32'b01110011100010001100110010011000;
		correct = 32'b01110011100010001100110010011000;
		#400 //1.8139834e-13 * 2.1676698e+31 = 2.1676698e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001111011111010110000000110;
		b = 32'b10110011010111111000101101000001;
		correct = 32'b10110011010111111000101101000001;
		#400 //5.7698927e-33 * -5.2047884e-08 = -5.2047884e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001110110101110101010000110;
		b = 32'b10001101000111111000110110010001;
		correct = 32'b11111001110110101110101010000110;
		#400 //-1.4208468e+35 * -4.916606e-31 = -1.4208468e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101000111011100101111000101000;
		b = 32'b00111001101100001000110110001111;
		correct = 32'b00111001101100001000110110001111;
		#400 //2.6464142e-14 * 0.00033674805 = 0.00033674805
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001001110011011011100101010;
		b = 32'b00011111001011101110001100011010;
		correct = 32'b01111001001110011011011100101010;
		#400 //6.026812e+34 * 3.7033787e-20 = 6.026812e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010110001111111110010111111;
		b = 32'b10001001011011000001001110100110;
		correct = 32'b01110010110001111111110010111111;
		#400 //7.922313e+30 * -2.8416705e-33 = 7.922313e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011001001111111010010111001111;
		b = 32'b00101000101100000100001110001010;
		correct = 32'b00101000101100000100001110001010;
		#400 //-9.907953e-24 * 1.9569216e-14 = 1.9569216e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101011100101110011111001010;
		b = 32'b11010010100000110100000000110000;
		correct = 32'b01010101011011101100110111001000;
		#400 //16692334000000.0 * -281858800000.0 = 16410474000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110000011101100110010010111;
		b = 32'b10101010101111010111111011100110;
		correct = 32'b01010110000011101100110010010111;
		#400 //39252340000000.0 * -3.3661198e-13 = 39252340000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000101100110001001000011011;
		b = 32'b01010100111000101011111100100000;
		correct = 32'b01010100111000101011111100100001;
		#400 //366736.84 * 7790953000000.0 = 7790954000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011100100011011101011111000;
		b = 32'b01010000111111101101001011001111;
		correct = 32'b01010000111111101101001011001111;
		#400 //-3.678751e-27 * 34201827000.0 = 34201827000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101001110011110000001011111;
		b = 32'b10000100011000001000100111011010;
		correct = 32'b01100101001110011110000001011111;
		#400 //5.4861045e+22 * -2.6394372e-36 = 5.4861045e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111101111000010000101010101;
		b = 32'b01010110100000100001000111110010;
		correct = 32'b01010110100000100001000111110010;
		#400 //96322.664 * 71506790000000.0 = 71506790000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011001011011111100110111100;
		b = 32'b01111100001011010001110000101011;
		correct = 32'b01111100001011010001110000101011;
		#400 //-2.103235e+26 * 3.5953547e+36 = 3.5953547e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110111100011100001010111010;
		b = 32'b11100100110010100101010111001110;
		correct = 32'b11100100110010100110010011101010;
		#400 //-8.7103454e+18 * -2.9859401e+22 = -2.9868111e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110000100100000111010001010;
		b = 32'b10010100011111011111111000011001;
		correct = 32'b11001110000100100000111010001010;
		#400 //-612606600.0 * -1.2823348e-26 = -612606600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010110011111101001100101111;
		b = 32'b01010110011010111011110000101001;
		correct = 32'b01010110011010111011110000101001;
		#400 //3.053713e-37 * 64798344000000.0 = 64798344000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010100100010001111001011001;
		b = 32'b01100110100101111000010101001011;
		correct = 32'b01100110100101111000010101001011;
		#400 //-3.933446e-18 * 3.5776808e+23 = 3.5776808e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010101000101001010001001110;
		b = 32'b11111000000000101110100110010011;
		correct = 32'b11111000000000101110100110010011;
		#400 //4.406721e-18 * -1.0620876e+34 = -1.0620876e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101001101010110110100111110;
		b = 32'b01011010100001010100111011110011;
		correct = 32'b01011010100001010100111011110011;
		#400 //-2.4011627e-21 * 1.8761489e+16 = 1.8761489e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000010100110001000000001011;
		b = 32'b11010000000011110111110001011111;
		correct = 32'b11010000000011110111110001011111;
		#400 //-2.727921e-24 * -9629171000.0 = -9629171000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010101100110000010111011111;
		b = 32'b10101011001111111010110011111101;
		correct = 32'b11000010101100110000010111011111;
		#400 //-89.51147 * -6.80969e-13 = -89.51147
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011100110100110011110001010;
		b = 32'b10000100011010111000110000000110;
		correct = 32'b10101011100110100110011110001010;
		#400 //-1.0971096e-12 * -2.7688413e-36 = -1.0971096e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101111001000001000111110000;
		b = 32'b00111110101000010110110010111101;
		correct = 32'b00111110101000010110110010111101;
		#400 //-3.956385e-16 * 0.31528273 = 0.31528273
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011110101011110001111010110;
		b = 32'b00101100100100011100111010100011;
		correct = 32'b11001011110101011110001111010110;
		#400 //-28034988.0 * 4.144089e-12 = -28034988.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111010110010011000010100000;
		b = 32'b11110011110101000010100011001011;
		correct = 32'b11110011110101000010100011001011;
		#400 //7.0177855e-25 * -3.361799e+31 = -3.361799e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111001110100001000001000101;
		b = 32'b11101001000011001101011001001001;
		correct = 32'b01111111001110100001000001000101;
		#400 //2.4732088e+38 * -1.0641347e+25 = 2.4732088e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001000000101011111110000000;
		b = 32'b01101000010101111100110011110101;
		correct = 32'b01101000010101111100110011110101;
		#400 //2300144000000000.0 * 4.0763583e+24 = 4.0763583e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000100011010001001000010111;
		b = 32'b11111000000100110100010010100100;
		correct = 32'b11111000000100110100010010100100;
		#400 //-5.5642566e-29 * -1.194781e+34 = -1.194781e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011110111001110010010010101;
		b = 32'b00000101110000010011101010001101;
		correct = 32'b01011011110111001110010010010101;
		#400 //1.2435165e+17 * 1.8171141e-35 = 1.2435165e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000000000001100001010100100;
		b = 32'b00010000010101111101111011111101;
		correct = 32'b10011000000000001100000111001100;
		#400 //-1.664188e-24 * 4.2573058e-29 = -1.6641455e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100000001101101111100110011;
		b = 32'b10110110100010011111000010010110;
		correct = 32'b10110110100010011111000010010110;
		#400 //1.0390151e-31 * -4.110926e-06 = -4.110926e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110000001001110111110101001;
		b = 32'b01010100010101111000111110001001;
		correct = 32'b01010100010101111000111110001001;
		#400 //2.5002515e-35 * 3703304400000.0 = 3703304400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010011101101100111110011001101;
		b = 32'b01110011000011010000110001110111;
		correct = 32'b01110011000011010000110001110111;
		#400 //1567555700000.0 * 1.1175029e+31 = 1.1175029e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110101010001001010111111000;
		b = 32'b00000101101100111101101110011001;
		correct = 32'b11000110101010001001010111111000;
		#400 //-21578.984 * 1.6913747e-35 = -21578.984
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000010111011000001100110001;
		b = 32'b10001001110000001110111110000011;
		correct = 32'b10111000010111011000001100110001;
		#400 //-5.2812687e-05 * -4.6447554e-33 = -5.2812687e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010010110011111010110011010001;
		b = 32'b10000001101111000000100111001101;
		correct = 32'b00010010110011111010110011010001;
		#400 //1.3106139e-27 * -6.9074357e-38 = 1.3106139e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100110110011111111101011001;
		b = 32'b11011011011010100101110001101000;
		correct = 32'b11111100110110011111111101011001;
		#400 //-9.05526e+36 * -6.5966746e+16 = -9.05526e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110001001000011001101000100;
		b = 32'b11000010000110101011001110000001;
		correct = 32'b11000010000110101011001110000001;
		#400 //-5.696841e-16 * -38.675297 = -38.675297
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101001001111010101100011100;
		b = 32'b11111111111101001010010011110101;
		correct = 32'b11111111111101001010010011110101;
		#400 //1.4542915e-16 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101010110111000100111101000;
		b = 32'b11011110011100010011100111000101;
		correct = 32'b11101101010110111000100111101000;
		#400 //-4.246496e+27 * -4.3455352e+18 = -4.246496e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100001101000111100011111100;
		b = 32'b10111110000110101110000101000110;
		correct = 32'b11010100001101000111100011111100;
		#400 //-3100495600000.0 * -0.15124997 = -3100495600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111101001001010110111111110;
		b = 32'b00000010111011100111011010001101;
		correct = 32'b11101111101001001010110111111110;
		#400 //-1.0193177e+29 * 3.5039002e-37 = -1.0193177e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110110001101100000000011011;
		b = 32'b01101000010111110101000110011011;
		correct = 32'b01101000010111110101000110011011;
		#400 //109264195000000.0 * 4.2183723e+24 = 4.2183723e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101001100101110110001100000;
		b = 32'b10100111111100110110000000111100;
		correct = 32'b00111101001100101110110001100000;
		#400 //0.043682456 * -6.7550386e-15 = 0.043682456
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010100001011000010011101000;
		b = 32'b01110111110101011100100001001011;
		correct = 32'b01110111110101011110100110101100;
		#400 //5.289239e+30 * 8.672044e+33 = 8.677333e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101110100011010011110111110;
		b = 32'b10001111101011111011100100010000;
		correct = 32'b01111101110100011010011110111110;
		#400 //3.4834952e+37 * -1.7327616e-29 = 3.4834952e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110111101010111100001001001;
		b = 32'b11010110111111101000011100101000;
		correct = 32'b11110110111101010111100001001001;
		#400 //-2.4893602e+33 * -139928220000000.0 = -2.4893602e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001111111110100001010110001;
		b = 32'b10110011101001001011111110111110;
		correct = 32'b01011001111111110100001010110001;
		#400 //8981181000000000.0 * -7.671723e-08 = 8981181000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001111011001011100001001100;
		b = 32'b01001000110001010100000101011111;
		correct = 32'b11010001111011001011100000011011;
		#400 //-127088030000.0 * 403978.97 = -127087630000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101000001111111111110010010001;
		b = 32'b11100011001101111000011011110001;
		correct = 32'b11100011001101111000011011110001;
		#400 //1.06573965e-14 * -3.3854777e+21 = -3.3854777e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011001110110001001010111010;
		b = 32'b10000010110011011110110010010110;
		correct = 32'b00001011001110110001001001010011;
		#400 //3.6028978e-32 * -3.0257836e-37 = 3.6028676e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010100101001100100010010100;
		b = 32'b10000101101111000101000010100010;
		correct = 32'b01111010100101001100100010010100;
		#400 //3.8626407e+35 * -1.7709055e-35 = 3.8626407e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100011011100010010111001101101;
		b = 32'b11111000011011001101010111000000;
		correct = 32'b11111000011011001101010111000000;
		#400 //-1.3074467e-17 * -1.9214335e+34 = -1.9214335e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101101010011101000110011110;
		b = 32'b10011011100100110001111100100011;
		correct = 32'b10011011100100110001111100100011;
		#400 //-1.5969685e-35 * -2.4339232e-22 = -2.4339232e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101000001101101110111110011;
		b = 32'b00000111101001110000000011101010;
		correct = 32'b11101101000001101101110111110011;
		#400 //-2.608707e+27 * 2.5127904e-34 = -2.608707e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100100010110100111111000010010;
		b = 32'b00100010011111110100010101010011;
		correct = 32'b10100100010010101000100110111101;
		#400 //-4.7378e-17 * 3.4595644e-18 = -4.3918437e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011111011111110100101001100;
		b = 32'b10100101110011011111011111001100;
		correct = 32'b10110011111011111110100101001100;
		#400 //-1.1171741e-07 * -3.5729745e-16 = -1.1171741e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011101111001101111001001000;
		b = 32'b01110001001000001010101111101110;
		correct = 32'b01110001001000001010101111101110;
		#400 //-4.767706e-27 * 7.956072e+29 = 7.956072e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001111111110100000010110010;
		b = 32'b00101111010001111010110001110100;
		correct = 32'b01000001111111110100000010110010;
		#400 //31.90659 * 1.8160212e-10 = 31.90659
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100100010101111000001011010;
		b = 32'b11010110011100111101000111100010;
		correct = 32'b11110100100010101111000001011010;
		#400 //-8.806297e+31 * -67020690000000.0 = -8.806297e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011011011001110011000110000;
		b = 32'b11101100000111000110011000100001;
		correct = 32'b11101100000111000110011000100001;
		#400 //2.9900879e-27 * -7.562989e+26 = -7.562989e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111111011110001010101000111;
		b = 32'b11100101011111101011010110011000;
		correct = 32'b11100101011111101011010110011000;
		#400 //-525749330000000.0 * -7.517693e+22 = -7.517693e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000101110010100110100000010;
		b = 32'b00011010010101001010001001110100;
		correct = 32'b01010000101110010100110100000010;
		#400 //24870654000.0 * 4.39718e-23 = 24870654000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001011110000111000011100000;
		b = 32'b10100110111010101100001111110001;
		correct = 32'b01001001011110000111000011100000;
		#400 //1017614.0 * -1.6290122e-15 = 1017614.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101000010110100001011110000;
		b = 32'b01011100000100100111101011111011;
		correct = 32'b01011101001011111110000110101111;
		#400 //6.271779e+17 * 1.6492226e+17 = 7.921002e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011101001100110101000000010;
		b = 32'b01110001010010000011011101000010;
		correct = 32'b01110001010010000011011101000010;
		#400 //-2.7530902e-22 * 9.914209e+29 = 9.914209e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111000100101100000110011010;
		b = 32'b00000000010001110011011011100001;
		correct = 32'b11101111000100101100000110011010;
		#400 //-4.541886e+28 * 6.540007e-39 = -4.541886e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001011011111011100010110101;
		b = 32'b01000111100001110001100100100011;
		correct = 32'b01001001100000000100110111101101;
		#400 //981899.3 * 69170.27 = 1051069.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000010000101000001000011100;
		b = 32'b10110011100010111000110100101000;
		correct = 32'b01110000010000101000001000011100;
		#400 //2.4078954e+29 * -6.498368e-08 = 2.4078954e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011111011101101010100001100;
		b = 32'b01101000000111001110110011110100;
		correct = 32'b01101000000111001110110011110100;
		#400 //3.9511475e-22 * 2.9642407e+24 = 2.9642407e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101010011001010111000010111;
		b = 32'b10111010110001101001101110110010;
		correct = 32'b01101101010011001010111000010111;
		#400 //3.9590877e+27 * -0.0015152602 = 3.9590877e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010111010100000101001101011111;
		b = 32'b11010001100001001100101110110101;
		correct = 32'b11010001100001001100101110110101;
		#400 //-6.7313654e-25 * -71294165000.0 = -71294165000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111010000111111000100010100;
		b = 32'b00001111001100011100101010101101;
		correct = 32'b01010111010000111111000100010100;
		#400 //215440190000000.0 * 8.765808e-30 = 215440190000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110111001011101111001011111;
		b = 32'b11100100111001110100001110010011;
		correct = 32'b11101110111001011101111001101101;
		#400 //-3.5570449e+28 * -3.4128537e+22 = -3.5570482e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000001001000110011110110000;
		b = 32'b10011000000101100110111101110011;
		correct = 32'b01110000001001000110011110110000;
		#400 //2.0352357e+29 * -1.9443313e-24 = 2.0352357e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101110001010001010000101111;
		b = 32'b00010001111101110011101101100000;
		correct = 32'b00010001111101110011101101100001;
		#400 //1.8533205e-35 * 3.9006321e-28 = 3.9006324e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110100001110010100101001110;
		b = 32'b10010000100100101010110111000011;
		correct = 32'b00100110100001110010100101001110;
		#400 //9.378702e-16 * -5.785457e-29 = 9.378702e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010011100010010001111110110;
		b = 32'b10101100101011101110111110111111;
		correct = 32'b10111010011100010010001111110110;
		#400 //-0.0009198779 * -4.9719946e-12 = -0.0009198779
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000100000010111011001110110;
		b = 32'b11100011100001101101111101001110;
		correct = 32'b11100011100001101101111101010000;
		#400 //-1138766300000000.0 * -4.975909e+21 = -4.97591e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		$display ("Done.");
		$finish;
	end

endmodule

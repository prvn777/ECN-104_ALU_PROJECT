`timescale 0.01 ns/1 ps
    `include "alu.v"


    module div_tb ();
        reg clock;
        reg [31:0] a, b;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] out;
        wire [49:0] pro;

        alu U1 (
                .clk(clock),
                .A(a),
                .B(b),
                .OPERATIONCODE(op),
                .O(out)
            );
       
        always
        #100 clock = ~clock; 
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clock, a, b, op, out);
            clock = 0;

    op = 3'b010;

		
		$display ("OPERATIONCODE: 010, Operation: DIV");
		
		a = 32'b00100001110010011001000010000101;
		b = 32'b10100111001000101111000001010010;
		correct = 32'b10111010000111100101011111100011;
		#400 //1.3658544e-18 * -2.2612294e-15 = -0.0006040318
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111110001000010101110010010;
		b = 32'b00011011010011000111011100001011;
		correct = 32'b01011011111101011001110101001111;
		#400 //2.338531e-05 * 1.6912949e-22 = 1.3826866e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001100011100001101000110000;
		b = 32'b11110000101011100010110001000110;
		correct = 32'b10101000010100001101110011001001;
		#400 //4999780000000000.0 * -4.3123132e+29 = -1.1594195e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010010011001100110101000111011;
		b = 32'b00010010100110111100001101011101;
		correct = 32'b00111111001111010101100010001110;
		#400 //7.2706142e-28 * 9.830036e-28 = 0.7396325
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001001000010001000101100001;
		b = 32'b10001101000111000001011010000111;
		correct = 32'b00111011100001000001010101110001;
		#400 //-1.9387842e-33 * -4.809833e-31 = 0.0040308763
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101001111010011011101010100;
		b = 32'b01010010101101011101100110100111;
		correct = 32'b00100010000001010010111101001000;
		#400 //7.04885e-07 * 390520340000.0 = 1.8049892e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100001111101001000101000001;
		b = 32'b01100111110011001001010010101010;
		correct = 32'b00110011111011100111011011101110;
		#400 //2.1455982e+17 * 1.9322103e+24 = 1.1104372e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110011000000000110010001101;
		b = 32'b10000101110010000011110001011110;
		correct = 32'b01011000000011110011100011110110;
		#400 //-1.1861057e-20 * -1.8830085e-35 = 629899200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011111000111011101100010110;
		b = 32'b10010011010101100001111001010101;
		correct = 32'b01100000000010000010001100101111;
		#400 //-1.0604542e-07 * -2.7025552e-27 = 3.9238944e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001101100001001000100111001111;
		b = 32'b10001101001010111101010000100111;
		correct = 32'b00111111110001010111011010000101;
		#400 //-8.168304e-31 * -5.2948812e-31 = 1.5426794
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		
		a = 32'b10100101010001111001010011010011;
		b = 32'b00010100010100010100100110000101;
		correct = 32'b11010000011101000010000010111001;
		#400 //-1.7310922e-16 * 1.0566303e-26 = -16383141000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100011011110100000110010100;
		b = 32'b10111101011100000111010010001000;
		correct = 32'b11010110011111101011100100110100;
		#400 //4110389600000.0 * -0.058704883 = -70017850000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101100110000100000011010011;
		b = 32'b01111010011010101001101010100011;
		correct = 32'b10100010101001100010001110000101;
		#400 //-1.3713751e+18 * 3.0453347e+35 = -4.5031998e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100111101110101010111110010;
		b = 32'b01001001100011001011000010110011;
		correct = 32'b10111010111000010000011010101110;
		#400 //-1978.6858 * 1152534.4 = -0.0017168128
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100000101110001011101011000;
		b = 32'b01100101110010100010010000010110;
		correct = 32'b00111101101111110101100100101111;
		#400 //1.1148562e+22 * 1.1932296e+23 = 0.09343182
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		$display ("Done.");
		$finish;
	end

endmodule

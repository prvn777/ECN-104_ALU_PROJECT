`timescale 0.01 ns/1 ps
    `include "alu.v"


    module add_tb ();
        reg clock;
        reg [31:0] a, b;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] out;
        wire [49:0] pro;

        alu U1 (
                .clk(clock),
                .A(a),
                .B(b),
                .OPERATIONCODE(op),
                .O(out)
            );
        
        always
        #100 clock = ~clock; 
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clock, a, b, op, out);
            clock = 0;

    op = 3'b000;

		
		$display ("OPERATIONCODE: 000, Operation: ADD");
	
		a = 32'b10110111001001011010001101000111;
		b = 32'b01000111110110100100000110001001;
		correct = 32'b01000111110110100100000110001001;
		#400 //-9.872782e-06 * 111747.07 = 111747.07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101110110101101010101101001;
		b = 32'b01011010010101101100100000000000;
		correct = 32'b01011010010101101100100000000000;
		#400 //458927400.0 * 1.5113887e+16 = 1.5113887e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		
		
		a = 32'b00110100101010100111001001001101;
		b = 32'b00101001110101011101111100111011;
		correct = 32'b00110100101010100111001001010000;
		#400 //3.1748132e-07 * 9.4978245e-14 = 3.174814e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000101001011000011111101001;
		b = 32'b11010001111101000111011110101110;
		correct = 32'b11010001111101000111011110101110;
		#400 //6.529043e-29 * -131247490000.0 = -131247490000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100000101100010100100010010;
		b = 32'b00100001110100100110101110001111;
		correct = 32'b00100001110100100110101110001111;
		#400 //-7.581164e-27 * 1.4258624e-18 = 1.4258624e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110010010111010101100100100;
		b = 32'b10011111010101000101000110010101;
		correct = 32'b10100110010010111010111001110101;
		#400 //-7.066171e-16 * -4.496023e-20 = -7.0666206e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001010111100111001010100110;
		b = 32'b00001110100011010010110110101100;
		correct = 32'b01010001010111100111001010100110;
		#400 //59712890000.0 * 3.4803164e-30 = 59712890000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001011011001011010100101001;
		b = 32'b01101111001011010010000100011000;
		correct = 32'b01101111001011010010000100011000;
		#400 //3.4445498e-09 * 5.3580915e+28 = 5.3580915e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000011110000110110001011100;
		b = 32'b10010101000011111000011001111101;
		correct = 32'b10111000011110000110110001011100;
		#400 //-5.9228725e-05 * -2.8984713e-26 = -5.9228725e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		
		a = 32'b11001111100100001110111111001100;
		b = 32'b11100011000111000010101010111100;
		correct = 32'b11100011000111000010101010111100;
		#400 //-4863269000.0 * -2.8807714e+21 = -2.8807714e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111000001010010010100010010100;
		b = 32'b01101011101101111010001100110000;
		correct = 32'b01111000001010010010100010010100;
		#400 //1.3723769e+34 * 4.440081e+26 = 1.3723769e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010010101110011010000010001;
		b = 32'b01100000111000011000100111101100;
		correct = 32'b01110010010101110011010000010001;
		#400 //4.2625422e+30 * 1.3001424e+20 = 4.2625422e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		
		a = 32'b11011000100000010111011001110110;
		b = 32'b11100011100001101101111101001110;
		correct = 32'b11100011100001101101111101010000;
		#400 //-1138766300000000.0 * -4.975909e+21 = -4.97591e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		$display ("Done.");
		$finish;
	end

endmodule

`timescale 0.01 ns/1 ps
    `include "alu.v"


    module sub_tb ();
        reg clock;
        reg [31:0] a, b;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] out;
        wire [49:0] pro;

        alu U1 (
                .clk(clock),
                .A(a),
                .B(b),
                .OPERATIONCODE(op),
                .O(out)
            );
        /* create a 10Mhz clock */
        always
        #100 clock = ~clock; // every 100 nanoseconds invert
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clock, a, b, op, out);
            clock = 0;

    op = 3'b001;

		/* Display the operation */
          $display ("OPERATIONCODE: 001, Operation: SUB");
		/* Test Cases!*/
		a = 32'b11111101110101110011001010100000;
		b = 32'b01000001010111010111101010010001;
		correct = 32'b11111101110101110011001010100000;
		#400 //-3.575586e+37 * 13.842423 = -3.575586e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011110110110011000101110111;
		b = 32'b00011110110111101110001001110110;
		correct = 32'b10110011110110110011000101110111;
		#400 //-1.020698e-07 * 2.3598826e-20 = -1.020698e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101100100000001111011110101110;
		b = 32'b01011101101110001111011100011101;
		correct = 32'b11011101101110001111011100011101;
		#400 //-3.6654768e-12 * 1.6660192e+18 = -1.6660192e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101100001110010001010101110;
		b = 32'b10110000100000110101110000100100;
		correct = 32'b11001101100001110010001010101110;
		#400 //-283399600.0 * -9.557692e-10 = -283399600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101110011100110110101101100;
		b = 32'b00001101100100110001001011001100;
		correct = 32'b11111101110011100110110101101100;
		#400 //-3.429864e+37 * 9.0641e-31 = -3.429864e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010010100110010100101010000;
		b = 32'b10001110111100100110010111011101;
		correct = 32'b10011010010100110010100101001110;
		#400 //-4.366715e-23 * -5.9755697e-30 = -4.3667143e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011010100111011101000101000;
		b = 32'b11011110110101101011010101010011;
		correct = 32'b01011110110101101011010101010011;
		#400 //1.1477753e-17 * -7.7356817e+18 = 7.7356817e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001011010111000011101111001;
		b = 32'b01011111110110110110000000111111;
		correct = 32'b01111001011010111000011101111001;
		#400 //7.643359e+34 * 3.1615408e+19 = 7.643359e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000001111000001001101110010;
		b = 32'b01100111001101110011011011010111;
		correct = 32'b11100111001101110011011011010111;
		#400 //12621564000.0 * 8.652047e+23 = -8.652047e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110100100101110001000011110;
		b = 32'b11000101110110011000110101011000;
		correct = 32'b01000101110110011000111110100100;
		#400 //0.2868814 * -6961.668 = 6961.955
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001010001101110011011100001;
		b = 32'b11001011000010011101010011000001;
		correct = 32'b11011001010001101110011011100001;
		#400 //-3499118700000000.0 * -9032897.0 = -3499118700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011010000000000011010100110;
		b = 32'b10101101111010100111011011001011;
		correct = 32'b00101101111010100111011011010001;
		#400 //1.0409749e-17 * -2.6655475e-11 = 2.6655485e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001011011000111100100010101;
		b = 32'b11100100100101010000000000110100;
		correct = 32'b11101001011011000010111010010101;
		#400 //-1.7867393e+25 * -2.1988636e+22 = -1.7845404e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100111010001101010001011101;
		b = 32'b11101010100000111000010010111111;
		correct = 32'b01101010100000111000010010111111;
		#400 //-5.2428552e+17 * -7.949808e+25 = 7.949808e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		$display ("Done.");
		$finish;
	end

endmodule

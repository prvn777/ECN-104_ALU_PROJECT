`timescale 0.01 ns/1 ps
    `include "alu.v"


    module div_tb ();
        reg clock;
        reg [31:0] a, b;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] out;
        wire [49:0] pro;

        alu U1 (
                .clk(clock),
                .A(a),
                .B(b),
                .OPERATIONCODE(op),
                .O(out)
            );
       
        always
        #100 clock = ~clock; 
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clock, a, b, op, out);
            clock = 0;

    op = 3'b010;

		
		$display ("OPERATIONCODE: 010, Operation: DIV");
		
		a = 32'b00100001110010011001000010000101;
		b = 32'b10100111001000101111000001010010;
		correct = 32'b10111010000111100101011111100011;
		#400 //1.3658544e-18 * -2.2612294e-15 = -0.0006040318
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111110001000010101110010010;
		b = 32'b00011011010011000111011100001011;
		correct = 32'b01011011111101011001110101001111;
		#400 //2.338531e-05 * 1.6912949e-22 = 1.3826866e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001100011100001101000110000;
		b = 32'b11110000101011100010110001000110;
		correct = 32'b10101000010100001101110011001001;
		#400 //4999780000000000.0 * -4.3123132e+29 = -1.1594195e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010010011001100110101000111011;
		b = 32'b00010010100110111100001101011101;
		correct = 32'b00111111001111010101100010001110;
		#400 //7.2706142e-28 * 9.830036e-28 = 0.7396325
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001001000010001000101100001;
		b = 32'b10001101000111000001011010000111;
		correct = 32'b00111011100001000001010101110001;
		#400 //-1.9387842e-33 * -4.809833e-31 = 0.0040308763
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101001111010011011101010100;
		b = 32'b01010010101101011101100110100111;
		correct = 32'b00100010000001010010111101001000;
		#400 //7.04885e-07 * 390520340000.0 = 1.8049892e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100001111101001000101000001;
		b = 32'b01100111110011001001010010101010;
		correct = 32'b00110011111011100111011011101110;
		#400 //2.1455982e+17 * 1.9322103e+24 = 1.1104372e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110011000000000110010001101;
		b = 32'b10000101110010000011110001011110;
		correct = 32'b01011000000011110011100011110110;
		#400 //-1.1861057e-20 * -1.8830085e-35 = 629899200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011111000111011101100010110;
		b = 32'b10010011010101100001111001010101;
		correct = 32'b01100000000010000010001100101111;
		#400 //-1.0604542e-07 * -2.7025552e-27 = 3.9238944e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001101100001001000100111001111;
		b = 32'b10001101001010111101010000100111;
		correct = 32'b00111111110001010111011010000101;
		#400 //-8.168304e-31 * -5.2948812e-31 = 1.5426794
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111011000101011100000010100;
		b = 32'b01101011101111011010011110100010;
		correct = 32'b10100011000110010000001111011010;
		#400 //-3803714600.0 * 4.585572e+26 = -8.294962e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000001100111001101010100100;
		b = 32'b00111110110000101111101011011000;
		correct = 32'b11010000111010111100111111110000;
		#400 //-12053025000.0 * 0.38082004 = -31650185000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101100101011110011111110011;
		b = 32'b11100100001101101011000111101000;
		correct = 32'b10000000110100100000111000000111;
		#400 //2.6004555e-16 * -1.3480508e+22 = -1.9290486e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111000110011111100010000100001;
		b = 32'b11001101111101010101011111001011;
		correct = 32'b01101010010110001100101001111100;
		#400 //-3.3711982e+34 * -514521440.0 = 6.5521046e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110001111101101100101100101;
		b = 32'b11010100101011111101000011110101;
		correct = 32'b11101001000010101111000111001010;
		#400 //6.3420524e+37 * -6041000000000.0 = -1.0498349e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100010111010100101111100001;
		b = 32'b10101100110010100101001111011110;
		correct = 32'b11100111000011000000000000011000;
		#400 //3801843200000.0 * -5.7504964e-12 = -6.6113304e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001110100100101000010011101011;
		b = 32'b10110001000001010011110000010000;
		correct = 32'b10011101000011001100001100111101;
		#400 //3.6119774e-30 * -1.9388189e-09 = -1.8629782e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110110100011101001110000001;
		b = 32'b01101110101110110110101010100100;
		correct = 32'b11001111100011110100111000011100;
		#400 //-1.3945342e+38 * 2.9001309e+28 = -4808521700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110011100001000101101001100;
		b = 32'b00111011001011010110110001101101;
		correct = 32'b10100010101100011000101001001010;
		#400 //-1.27343e-20 * 0.0026462332 = -4.8122365e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010110010001001100100010101;
		b = 32'b01101011100011011010001010101010;
		correct = 32'b00011110101101010100100101000011;
		#400 //6573194.5 * 3.424534e+26 = 1.919442e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011011010011111110011100000;
		b = 32'b00101001011111111101010001111111;
		correct = 32'b00100001011010100010010010101010;
		#400 //4.506441e-32 * 5.6805685e-14 = 7.933081e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011110101100010110100110011;
		b = 32'b11010010100001101110110010010011;
		correct = 32'b11100000110010110010111101110001;
		#400 //3.393763e+31 * -289747340000.0 = -1.1712836e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110001010000110100110010111;
		b = 32'b11011010010100111110100001010100;
		correct = 32'b11001011010010110111010001101001;
		#400 //1.9882634e+23 * -1.4911667e+16 = -13333609.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100001111011101001111100010;
		b = 32'b01000101000001000000001111101101;
		correct = 32'b01001110101110000000110111001110;
		#400 //3261214500000.0 * 2112.2454 = 1543956200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110101101010000111000000010011;
		b = 32'b01011011010010101000101100011101;
		correct = 32'b11011001110101001110010010011100;
		#400 //-4.2704053e+32 * 5.70109e+16 = -7490506700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010010100010010011001000001;
		b = 32'b10000011111000111111011101001100;
		correct = 32'b01100101111010101101111010010101;
		#400 //-1.8576201e-13 * -1.33986375e-36 = 1.3864246e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110001000001000101111000111;
		b = 32'b01000101000111100011011010001000;
		correct = 32'b01000000100000011110001100110010;
		#400 //10274.944 * 2531.4082 = 4.058984
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011110101111001000010110001;
		b = 32'b01101010101011100110100101101000;
		correct = 32'b00110000100111100011001111001100;
		#400 //1.2135242e+17 * 1.0542543e+26 = 1.1510735e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101000110000101100111100000;
		b = 32'b00100100010101001101010110011001;
		correct = 32'b01110000001101110011111111111001;
		#400 //10469486000000.0 * 4.6151096e-17 = 2.2685238e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001011101111000011110001101;
		b = 32'b00000110101101001001000011001110;
		correct = 32'b10111010001011110111100000110110;
		#400 //-4.5463988e-38 * 6.7921246e-35 = -0.0006693633
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010010110110001110011011110;
		b = 32'b10011100011011101111101011001101;
		correct = 32'b01101101011010101011011111011000;
		#400 //-3589943.5 * -7.9071747e-22 = 4.540109e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011100111110110100001110111;
		b = 32'b10100010101110001010110001110001;
		correct = 32'b11100000010111001111100111100110;
		#400 //318.81613 * -5.005588e-18 = -6.3692043e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011011011000110001110001100;
		b = 32'b10110100000000100111100011001110;
		correct = 32'b00110110111001111110100100001000;
		#400 //-8.398219e-13 * -1.2151142e-07 = 6.911465e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111001101001110000010010110011;
		b = 32'b00100001101000000000010111100001;
		correct = 32'b11010111100001011001100001110011;
		#400 //-0.00031856223 * 1.0843578e-18 = -293779620000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110000011101110101111101111;
		b = 32'b10010100001010100010110000111011;
		correct = 32'b01011001010101110000000100101111;
		#400 //-3.2496613e-11 * -8.5915296e-27 = 3782401300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111111000101101000110010100;
		b = 32'b10110111100001000111011101011010;
		correct = 32'b00010111110110110010101111011000;
		#400 //-2.2366047e-29 * -1.5791204e-05 = 1.4163611e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100000101110010110011011110;
		b = 32'b00101100101111001011011010111000;
		correct = 32'b11101110110011010001001110111101;
		#400 //-1.7020821e+17 * 5.3635672e-12 = -3.1734145e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110001100011000100011001001;
		b = 32'b01000001100000110001101110111001;
		correct = 32'b10100100001011010101001101001011;
		#400 //-6.159459e-16 * 16.388536 = -3.7583947e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010011000011010100001111001;
		b = 32'b00011010000100110110101111111110;
		correct = 32'b11001111110000111110110111011101;
		#400 //-2.0042465e-13 * 3.0486123e-23 = -6574291500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111110110101000110100000000;
		b = 32'b01001010010101000111011011100010;
		correct = 32'b11011101000000111010101010110010;
		#400 //-2.0641538e+24 * 3481016.5 = -5.9297445e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110110001111011110101011001100;
		b = 32'b01001110111010010100111110011000;
		correct = 32'b01100110110100000110001011100100;
		#400 //9.629945e+32 * 1957153800.0 = 4.9203822e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001100100011101010000010001;
		b = 32'b10000000000010100000000101100111;
		correct = 32'b01001010011010010011001010011011;
		#400 //-3.5106907e-33 * -9.18858e-40 = 3820710.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011101010011101100100011000;
		b = 32'b11010010101110000110010100001010;
		correct = 32'b11011000011010111100110111110011;
		#400 //4.1066732e+26 * -395984570000.0 = -1037079100000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101010000110001110011101100000;
		b = 32'b10011010011101100000000001001010;
		correct = 32'b11001111000111110001111001100010;
		#400 //1.3580586e-13 * -5.087184e-23 = -2669568500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110100111101010101010100000;
		b = 32'b01001111100111010101000111100010;
		correct = 32'b01000110100000010001100001111110;
		#400 //87227830000000.0 * 5278778400.0 = 16524.246
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101111010000000000010110111001;
		b = 32'b10001100110101110010110010001110;
		correct = 32'b01100001111001000111010010100101;
		#400 //-1.7464331e-10 * -3.315281e-31 = 5.2678285e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100000111110000110011110111110;
		b = 32'b01011101001010001101000111110000;
		correct = 32'b11000011001111000101011101111110;
		#400 //-1.4319587e+20 * 7.60298e+17 = -188.34177
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011111001110111111100011001;
		b = 32'b11110101011011010001101100000101;
		correct = 32'b00000101111110011111000110100111;
		#400 //-0.007064712 * -3.0056699e+32 = 2.3504617e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110010100100110110011010010;
		b = 32'b00010010001010100001110110011011;
		correct = 32'b00110011100111100101010001111011;
		#400 //3.957656e-35 * 5.3679033e-28 = 7.372815e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011111000111110011111111000;
		b = 32'b11100000011000110101011100100111;
		correct = 32'b10000011000000000101000110001001;
		#400 //2.4709632e-17 * -6.552642e+19 = -3.7709417e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100011110110110001101100101;
		b = 32'b01110010100110001101001011000011;
		correct = 32'b00010001010100101000111000010000;
		#400 //1005.55304 * 6.053954e+30 = 1.6609855e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011100110011000100011001101;
		b = 32'b00111100111000011000110000111001;
		correct = 32'b00011110001011100100001110000111;
		#400 //2.5400132e-22 * 0.027532684 = 9.225448e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110010010100111000000111011;
		b = 32'b01101111011101101001110110111111;
		correct = 32'b10101110010100100010010000101000;
		#400 //-3.646806e+18 * 7.6324016e+28 = -4.7780585e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010001101100110001011001000;
		b = 32'b00001001111101001100000001010011;
		correct = 32'b11110111101111101100010010101111;
		#400 //-45.596466 * 5.8921724e-33 = -7.7384814e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100111010111101001110111001;
		b = 32'b11100000001100010001011110111000;
		correct = 32'b00100100001010100111001111001110;
		#400 //-1886.6163 * -5.104348e+19 = 3.6960964e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101101011001101110100100101;
		b = 32'b10001111001000011001011000001110;
		correct = 32'b01001110000010001110111100000000;
		#400 //-4.575668e-21 * -7.966812e-30 = 574341100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000000000000001000001110000;
		b = 32'b11101011110001101100100110000000;
		correct = 32'b00011011101001001110110000011111;
		#400 //-131137.75 * -4.8063774e+26 = 2.7284114e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000111001110001101101111111;
		b = 32'b10000111100111000111100000011001;
		correct = 32'b11000000101111010000111011011100;
		#400 //1.3909271e-33 * -2.3542858e-34 = -5.908064
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000100110110000101111101001;
		b = 32'b10111110101100001111100100110001;
		correct = 32'b01001001011000000100100000100011;
		#400 //-317535.28 * -0.34565118 = 918658.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101110001101011101111111001;
		b = 32'b01100000111001011011100101101000;
		correct = 32'b10100100010111010111011100100101;
		#400 //-6359.4966 * 1.3242701e+20 = -4.8022655e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111001001110001100010010010;
		b = 32'b10110110000010110011111001001000;
		correct = 32'b01101000100110011001101010001101;
		#400 //-1.2040534e+19 * -2.0748867e-06 = 5.802984e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100001110111100000011000000;
		b = 32'b01010011110101110000000100110101;
		correct = 32'b10100111110111111000110101010101;
		#400 //-0.011459529 * 1846876400000.0 = -6.2048166e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111111001100000110011111101;
		b = 32'b01000001000111111100010111000010;
		correct = 32'b00111110001110000100110101111011;
		#400 //1.7972714 * 9.985781 = 0.17998306
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110010101111010010110100010;
		b = 32'b00100010100101011100111011110100;
		correct = 32'b01010011001110000100000100001110;
		#400 //3.2133908e-06 * 4.060565e-18 = 791365400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100011000000011110011011100;
		b = 32'b11010100010110000011010100001011;
		correct = 32'b11010111100001001100000100011000;
		#400 //1.0843471e+27 * -3714411400000.0 = -291929730000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110000100010111010100001110;
		b = 32'b01111010111111111000101110110010;
		correct = 32'b10111010100100011011011101000001;
		#400 //-7.3755586e+32 * 6.6343453e+35 = -0.0011117236
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001001000001000010010000000;
		b = 32'b00101011111011110110011101101001;
		correct = 32'b10100100101010111010010100100001;
		#400 //-1.2662604e-28 * 1.7010673e-12 = -7.443917e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000000010010101010100001100;
		b = 32'b00011000101000000110110110001111;
		correct = 32'b00101110110110110010010100111000;
		#400 //4.132691e-34 * 4.1469657e-24 = 9.9655784e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010110011101000110110010110;
		b = 32'b01110100011100110110100001101101;
		correct = 32'b00101101110110010011110100010011;
		#400 //1.9051158e+21 * 7.7139047e+31 = 2.4697166e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001011110101000011010111010;
		b = 32'b10101011110000010100011001110010;
		correct = 32'b01111101001001011110101001100100;
		#400 //-1.892923e+25 * -1.3733027e-12 = 1.3783728e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101100101111110001011110110100;
		b = 32'b01100110101001100010101101100110;
		correct = 32'b10000101100100110011001010111100;
		#400 //-5.431178e-12 * 3.923567e+23 = -1.384245e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111101010100101111110110110;
		b = 32'b00010101110110000001010001110101;
		correct = 32'b01111001010010011101100110010100;
		#400 //5716798500.0 * 8.727398e-26 = 6.550404e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100101101111001010100011001;
		b = 32'b11101000111010101111111000010110;
		correct = 32'b10001011010001111111111001111000;
		#400 //3.419489e-07 * -8.8777665e+24 = -3.8517447e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111000101101001110001011001110;
		b = 32'b10010110110010110101110111001001;
		correct = 32'b11100001011000111011001110010000;
		#400 //8.6253145e-05 * -3.2855606e-25 = -2.6252186e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000001100011001100101100010;
		b = 32'b10011110101010001011010100010111;
		correct = 32'b11101001000001101011111100001100;
		#400 //181861.53 * -1.7862589e-20 = -1.0181141e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001111111011110011101001111;
		b = 32'b10000011000001001000001111111011;
		correct = 32'b01000110011101010100000001101011;
		#400 //-6.1125056e-33 * -3.894282e-37 = 15696.1045
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101001010000110110111100011;
		b = 32'b10010101111001110000001101110000;
		correct = 32'b01100110101110101010010110001100;
		#400 //-0.04112042 * -9.330558e-26 = 4.40707e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000100110010011100101011001;
		b = 32'b11000101100101000101001111011110;
		correct = 32'b11000010100001000011100110110010;
		#400 //313802.78 * -4746.4834 = -66.112686
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111111101001011010111001111;
		b = 32'b10110111000111000000111000001000;
		correct = 32'b01011000010010001011011110100011;
		#400 //-8211111400.0 * -9.3015915e-06 = 882764160000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100010000111101100010011001;
		b = 32'b01110110001101010111110011001111;
		correct = 32'b00010101100010100010000001111000;
		#400 //51339876.0 * 9.202511e+32 = 5.578898e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010000001010000101111000101;
		b = 32'b11011000010001101001110010101110;
		correct = 32'b00010001001010110111110100101100;
		#400 //-1.1816856e-13 * -873504950000000.0 = 1.3528093e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100010100110101111110011010;
		b = 32'b11110001101110000101010110100100;
		correct = 32'b11001010000100101100011010001010;
		#400 //4.3900547e+36 * -1.8255608e+30 = -2404770.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001110101000100001110111001;
		b = 32'b01010111001101110110000011111111;
		correct = 32'b00010010000101000010100110010101;
		#400 //9.426439e-14 * 201627220000000.0 = 4.675182e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110111001000111000101001001010;
		b = 32'b01010011010010110111111011111000;
		correct = 32'b01100011010011011011110000111000;
		#400 //3.316989e+33 * 874008540000.0 = 3.795145e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001000111101110110010010011;
		b = 32'b11101001001101100101011011111011;
		correct = 32'b00011111010111110010000000000101;
		#400 //-650953.2 * -1.3777203e+25 = 4.7248573e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010000111110110100001000011;
		b = 32'b10111001000100101100111110110010;
		correct = 32'b00010000100010101111101101100101;
		#400 //-7.675181e-33 * -0.00014001018 = 5.481874e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111010111111110101110000001;
		b = 32'b11111111011100011001000011000111;
		correct = 32'b00001111011011010100110011001101;
		#400 //-3756753200.0 * -3.2109567e+38 = 1.16997935e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110011111001100111101001101;
		b = 32'b01010101010000001101100110101010;
		correct = 32'b00100000101001111100101111111010;
		#400 //3.7671591e-06 * 13252568000000.0 = 2.842588e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010111100000110010000110010;
		b = 32'b01100100010010011111101010000100;
		correct = 32'b01000110000110000101011111100111;
		#400 //1.4530768e+26 * 1.4903388e+22 = 9749.976
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000001000011001000110010110;
		b = 32'b00011000100100110101000010000111;
		correct = 32'b11101111000011000110001010100000;
		#400 //-165446.34 * 3.807992e-24 = -4.344713e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011010000000011001011010000;
		b = 32'b10111001010110001001010000011000;
		correct = 32'b01111001011000110010111010101111;
		#400 //-1.5227533e+31 * -0.00020654534 = 7.372489e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101000010101010111010001100111;
		b = 32'b01100100110000111101010110000101;
		correct = 32'b00000011000010111000010001100001;
		#400 //1.1849116e-14 * 2.8900006e+22 = 4.100039e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011101110111000111000100001;
		b = 32'b01100001101111001110000001010101;
		correct = 32'b00111001011111100011010110011011;
		#400 //1.0558419e+17 * 4.355191e+20 = 0.00024243297
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111000100001011100111011101100;
		b = 32'b11100000110100111010101001010010;
		correct = 32'b11010111001000011101010111010111;
		#400 //2.1711636e+34 * -1.2201675e+20 = -177939800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110111100101000010100001111000;
		b = 32'b01101101101111000100001000101000;
		correct = 32'b11001001010010010111100001100001;
		#400 //-6.010006e+33 * 7.282895e+27 = -825222.06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101110100000011101110011011;
		b = 32'b01000000110101000110010010011011;
		correct = 32'b01010100011110101111110001011000;
		#400 //28619303000000.0 * 6.637281 = 4311901800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111011001010110010011001001;
		b = 32'b11110010001000100011111000101111;
		correct = 32'b10100100101101001111101001011101;
		#400 //252221030000000.0 * -3.2135518e+30 = -7.848669e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111010100100101110111100000;
		b = 32'b01011000110000001100110100010101;
		correct = 32'b00110110000010111010100101101000;
		#400 //3529367600.0 * 1695896400000000.0 = 2.0811221e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001110010001000110011111101;
		b = 32'b10000011100111110000111110011010;
		correct = 32'b11101101101000010110001101000110;
		#400 //5.8367946e-09 * -9.348762e-37 = -6.2433876e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111001001100001101100111010011;
		b = 32'b10000100010111011011100111100100;
		correct = 32'b01110100010011000011000000100011;
		#400 //-0.00016865814 * -2.6063782e-36 = 6.470977e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010011011010001110000110100;
		b = 32'b00100001001001001100100010011001;
		correct = 32'b01101000101110000010111001111100;
		#400 //3884813.0 * 5.583085e-19 = 6.9581833e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010010010101001101100100011000;
		b = 32'b00110011101011000001110011101011;
		correct = 32'b11011110000111100100101101101001;
		#400 //-228543820000.0 * 8.014634e-08 = -2.8515815e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011001110110000111111000110;
		b = 32'b10000110100101010010110101111111;
		correct = 32'b01010100001000001000000101111011;
		#400 //-1.5473374e-22 * -5.611442e-35 = 2757468400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011010011111011110000101001;
		b = 32'b11010101101011110010110011110010;
		correct = 32'b01010101000101111100101010000001;
		#400 //-2.511362e+26 * -24075947000000.0 = 10431000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011011101110101110001100011;
		b = 32'b00100001000110010011101111001010;
		correct = 32'b01001001110011101010000010000101;
		#400 //8.788024e-13 * 5.1917547e-19 = 1692688.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101100111111011111101011110;
		b = 32'b11011010011000001101011100001010;
		correct = 32'b10111010101101011110001011110100;
		#400 //21955533000000.0 * -1.5821708e+16 = -0.0013876841
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001101010011000101000100010001;
		b = 32'b00010011111110110101101010111111;
		correct = 32'b10111000110100000001011111000100;
		#400 //-6.2959934e-31 * 6.345079e-27 = -9.9226396e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101001000100100010010101111;
		b = 32'b00110110001000010110101001001100;
		correct = 32'b01110110100000001010110100101101;
		#400 //3.1387253e+27 * 2.4052742e-06 = 1.3049344e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101111111110010010011001010;
		b = 32'b00110000000011110101110100101100;
		correct = 32'b01110101011000111100110011110100;
		#400 //1.5061026e+23 * 5.21555e-10 = 2.8877156e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111100001100001000101001101;
		b = 32'b01100110000010001010101111110010;
		correct = 32'b10111000111110110001111101001110;
		#400 //-1.9321175e+19 * 1.6135342e+23 = -0.000119744436
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010111001011011011000110010;
		b = 32'b01111001111000000000110001111111;
		correct = 32'b01000000100000110011110000111000;
		#400 //5.9636567e+35 * 1.4541599e+35 = 4.101101
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110111001001001011000101010;
		b = 32'b00100111011011111110100111110111;
		correct = 32'b01011110111100111110100111000101;
		#400 //29259.082 * 3.3294745e-15 = 8.787898e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001011100010101110111110110;
		b = 32'b01110011010001001000011100011101;
		correct = 32'b00100101100111010011010001000010;
		#400 //4246173800000000.0 * 1.5570535e+31 = 2.727057e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101101110001001100000011010;
		b = 32'b00111100010011001101110010101100;
		correct = 32'b01010000111001101010110001000000;
		#400 //387122000.0 * 0.012503784 = 30960386000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101000001110000111110011110;
		b = 32'b00010110001000010110110011010000;
		correct = 32'b01101110010101100011000010011110;
		#400 //2160.976 * 1.3039812e-25 = 1.6572142e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011110100001010001110111001;
		b = 32'b10111110010010000100001010011010;
		correct = 32'b11011101000001010101101100011000;
		#400 //1.1745362e+17 * -0.19556656 = -6.005813e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111011001000111001010101010;
		b = 32'b11101110001101101010011001001000;
		correct = 32'b01010000101000000001100001100101;
		#400 //-3.0365935e+38 * -1.4131823e+28 = 21487626000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111000100100010110100100001;
		b = 32'b01010011010111001100101111000110;
		correct = 32'b01101011001010010111101110011011;
		#400 //1.943016e+38 * 948311560000.0 = 2.0489217e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001001010101011111110010010;
		b = 32'b00001100000111100001101010100101;
		correct = 32'b11100100100010100011110010011000;
		#400 //-2.484715e-09 * 1.2179895e-31 = -2.0400135e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111110101010000101010000001;
		b = 32'b11011101010011111011001100101001;
		correct = 32'b10101010000000110100101010101001;
		#400 //109077.01 * -9.3539694e+17 = -1.166104e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001101001111100111101010111;
		b = 32'b11001010000011011000111100100000;
		correct = 32'b10110111000101111011110010000111;
		#400 //20.97624 * -2319304.0 = -9.044196e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010010010111001110110000110011;
		b = 32'b11011010011100011111100000110111;
		correct = 32'b00110111011010011011101110010001;
		#400 //-237213900000.0 * -1.7027096e+16 = 1.3931553e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000101111101011101111001110;
		b = 32'b00110000110100000000001110100000;
		correct = 32'b10111111011010101011101110101011;
		#400 //-1.3877697e-09 * 1.5135022e-09 = -0.9169261
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010011100101011101000101011;
		b = 32'b01111010000010011001011011000011;
		correct = 32'b10000111111000011100111110011011;
		#400 //-60.681805 * 1.7860062e+35 = -3.3976257e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111000101110000001000000011;
		b = 32'b01101110101001101000111111101011;
		correct = 32'b01001111111010000001011111110101;
		#400 //2.0072387e+38 * 2.577425e+28 = 7787768300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111111000011101101110110101;
		b = 32'b11100100000011000011110011100011;
		correct = 32'b11111111111000011101101110110101;
		#400 //nan * -1.0347726e+22 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111010110111001010011010000;
		b = 32'b11001001110111101001011001110111;
		correct = 32'b11100100111111001000101011010001;
		#400 //6.795712e+28 * -1823438.9 = -3.7268658e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010011000101011110101110100;
		b = 32'b01001100000100100000000010000001;
		correct = 32'b10011101110001101100100001111010;
		#400 //-2.0138562e-13 * 38273540.0 = -5.261745e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011010011000101111011111011;
		b = 32'b11011001011111010010111011100100;
		correct = 32'b11100001010011101010010100010000;
		#400 //1.061155e+36 * -4454045400000000.0 = -2.382452e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110000000000001100000111101;
		b = 32'b11111001000110110110110000101001;
		correct = 32'b00011100010100101111110011011011;
		#400 //-35210398000000.0 * -5.0437485e+34 = 6.980998e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001000110110100011101001001110;
		b = 32'b10001101101000011101000101111100;
		correct = 32'b00111010101011001001111011011000;
		#400 //-1.3134105e-33 * -9.972823e-31 = 0.0013169898
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100110011000011111100011011;
		b = 32'b11111000100011110001011111100101;
		correct = 32'b00001011101101101011001111101010;
		#400 //-1633.972 * -2.3218222e+34 = 7.0374555e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001110000100001010010001111;
		b = 32'b11010010101100100001101101000100;
		correct = 32'b01001110100010110111101011011011;
		#400 //-4.4751872e+20 * -382480800000.0 = 1170042200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011001011011001110100111000;
		b = 32'b01110101010011011000111101011011;
		correct = 32'b00101101010110000011011100100000;
		#400 //3.2026155e+21 * 2.6057823e+32 = 1.2290419e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010101110000111110101001010;
		b = 32'b00101111100110000100011110001011;
		correct = 32'b11010010100110110001001100001011;
		#400 //-92.244705 * 2.7699473e-10 = -333019700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001000001111000111101110000;
		b = 32'b11111000101010101001110111010100;
		correct = 32'b10100111110010110110011001110101;
		#400 //1.5629039e+20 * -2.7684113e+34 = -5.6454903e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001000110110111011011111100;
		b = 32'b01000111111001110110100001011100;
		correct = 32'b00100000101010111111110010001001;
		#400 //3.4520116e-14 * 118480.72 = 2.913564e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101110010101110000000100111;
		b = 32'b11110000000111011011111110011001;
		correct = 32'b00010101001001001001110111110101;
		#400 //-6492.019 * -1.952831e+29 = 3.3244142e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100011000011101000001101010000;
		b = 32'b00010111010011111100110011110110;
		correct = 32'b11001011001011111001000110011111;
		#400 //-7.725642e-18 * 6.7144004e-25 = -11506079.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111010110010101100110100000;
		b = 32'b01001110000000111011110011011100;
		correct = 32'b00111000110100110010111011101111;
		#400 //55641.625 * 552548100.0 = 0.00010070006
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001101011010100110101000001;
		b = 32'b01101110001001100100101000110101;
		correct = 32'b00011011000001010110010110111000;
		#400 //1419688.1 * 1.2866056e+28 = 1.1034369e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010111001011111110010111101;
		b = 32'b01000000110011110010011111010110;
		correct = 32'b01011001100011100001101110000110;
		#400 //3.236783e+16 * 6.473613 = 4999963600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000011111001110000011011111;
		b = 32'b10100111001110110011010100111110;
		correct = 32'b11110000101011001110011010100100;
		#400 //1112171000000000.0 * -2.5980326e-15 = -4.28082e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110111111111000011101101001;
		b = 32'b01100110101000001100100001011110;
		correct = 32'b11000111110010110110110110010100;
		#400 //-3.954119e+28 * 3.7963738e+23 = -104155.16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000001101110000101110111000;
		b = 32'b00110010111111010010010110100011;
		correct = 32'b10111100101110010001101111010101;
		#400 //-6.6591666e-10 * 2.9470192e-08 = -0.02259628
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110001000010010000110101111;
		b = 32'b01110010101011001110111011001100;
		correct = 32'b00000010111011101000011110110111;
		#400 //2.4010476e-06 * 6.850574e+30 = 3.5048853e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010101000110100100111000110;
		b = 32'b00101000011111000100110011101110;
		correct = 32'b10101001101001011010111010110111;
		#400 //-1.0304933e-27 * 1.4005492e-14 = -7.35778e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011010010101000111100001101;
		b = 32'b00110101110010100001011010111111;
		correct = 32'b10001101000000000100110000110011;
		#400 //-5.952668e-37 * 1.5056793e-06 = -3.9534767e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001101001101010000001001110;
		b = 32'b10010111111101010110010101110110;
		correct = 32'b11111001001011011101001110000000;
		#400 //89456755000.0 * -1.5858366e-24 = -5.640982e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000000000011100111100111000;
		b = 32'b01001100100110010000001000100110;
		correct = 32'b11100010110110010010111110000011;
		#400 //-1.6069631e+29 * 80220460.0 = -2.0031835e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010100010100101111000010010;
		b = 32'b00010011000010010010101110000011;
		correct = 32'b01001111000000010001111000010001;
		#400 //3.7504576e-18 * 1.7313284e-27 = 2166231300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101111010111000101111101011;
		b = 32'b01101100111010101010010001111110;
		correct = 32'b00001000100000000111111000111111;
		#400 //1.7549586e-06 * 2.2693235e+27 = 7.7334e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000100101010011011100011000;
		b = 32'b10110011100110010101001110011000;
		correct = 32'b11111100011110010010001010110100;
		#400 //3.6943897e+29 * -7.139823e-08 = -5.174343e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000110111001100111001011011010;
		b = 32'b00011000100101100001101000111000;
		correct = 32'b10101101110001001000001111101101;
		#400 //-8.6685143e-35 * 3.8800565e-24 = -2.2341207e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111010111011101101101100111;
		b = 32'b11000000110111100011110111010101;
		correct = 32'b11001101111111111000111010011110;
		#400 //3722143500.0 * -6.945048 = -535942080.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111111100110010100001011101;
		b = 32'b10011011001011001110110000000000;
		correct = 32'b11111100001100111111110101100111;
		#400 //534709370000000.0 * -1.4303762e-22 = -3.738243e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110010110001110111101001000;
		b = 32'b00001000011010001100101011100011;
		correct = 32'b11100101011011101000111110110000;
		#400 //-4.932524e-11 * 7.0053453e-34 = -7.041086e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110100011000100011000111111001;
		b = 32'b11100110111010001100010001000101;
		correct = 32'b00001100111110001100010111001001;
		#400 //-2.106607e-07 * -5.4960478e+23 = 3.8329488e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110001111110000110010100110;
		b = 32'b01100011111011110100011111101111;
		correct = 32'b10000001110011000110010111111101;
		#400 //-6.628358e-16 * 8.8279104e+21 = -7.508411e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011110110101100100100111010100;
		b = 32'b00100011010001000000101110110001;
		correct = 32'b00111011000010111110100100101101;
		#400 //2.2688666e-20 * 1.0627657e-17 = 0.00213487
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001000110101110011011111111;
		b = 32'b11000011001111000011100111111011;
		correct = 32'b00001101010100101010110101010001;
		#400 //-1.2219639e-28 * -188.22649 = 6.491987e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111100000100100011001111101;
		b = 32'b11001000011101100001000010011010;
		correct = 32'b00000110100001111000100100001101;
		#400 //-1.2846141e-29 * -251970.4 = 5.0982734e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001000111101100010110110011;
		b = 32'b11001011111101101110011111010100;
		correct = 32'b10011100101001001001111011010100;
		#400 //3.5254524e-14 * -32362408.0 = -1.0893666e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001110010101011011000001100;
		b = 32'b10101100011101011100001101001000;
		correct = 32'b11101100110100110010011110101110;
		#400 //7132263500000000.0 * -3.4924997e-12 = -2.0421658e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000101111011011101111110001;
		b = 32'b01001111110110010010110110101001;
		correct = 32'b01000000010111111010011001100111;
		#400 //25465686000.0 * 7287296500.0 = 3.4945314
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001110000001110010100001111;
		b = 32'b11110000100001110010010101110010;
		correct = 32'b10110000101101101011000111100010;
		#400 //4.4478503e+20 * -3.3460596e+29 = -1.32928e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110001000010011110111011001;
		b = 32'b01101011101000010010101001111011;
		correct = 32'b10010010000000000000111101100010;
		#400 //-0.1574625 * 3.8967533e+26 = -4.040864e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101100110011001001011011100001;
		b = 32'b11010000010101110110010011100111;
		correct = 32'b00011011111100110010100010000111;
		#400 //-5.8147796e-12 * -14454857000.0 = 4.0227168e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100101111111010010001000101;
		b = 32'b10000101111001000000011111000011;
		correct = 32'b11101110010101110010010111100100;
		#400 //3.5696044e-07 * -2.1443868e-35 = -1.6646271e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111011110111010110011100101;
		b = 32'b00011000011011001101011010000100;
		correct = 32'b11111110100010000000010011011001;
		#400 //-276720000000000.0 * 3.0610588e-24 = -9.040009e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111100100111110101111110011;
		b = 32'b01100010111101011100101000000110;
		correct = 32'b00100100000110100001000100011010;
		#400 //75735.9 * 2.2670048e+21 = 3.3407912e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011111001000100100011010001;
		b = 32'b10110000110110010100100110011111;
		correct = 32'b01011010100001100111101001100001;
		#400 //-29921698.0 * -1.5809752e-09 = 1.8926102e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000100010001101000110101000;
		b = 32'b11010001001010010100100000010011;
		correct = 32'b11001110110011101110100001100000;
		#400 //7.887077e+19 * -45441167000.0 = -1735667700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010010000010110100110000000;
		b = 32'b00101000110000100110010011001100;
		correct = 32'b01101000111111101011010100010000;
		#400 //207674670000.0 * 2.158204e-14 = 9.622569e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010010001010101001111000001110;
		b = 32'b00110110000100011110110110010100;
		correct = 32'b00011011100101011010011111111001;
		#400 //5.383736e-28 * 2.1744972e-06 = 2.4758532e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000001001110010010001011001011;
		b = 32'b00001010000100110101011010010100;
		correct = 32'b00110110101000001101011000110101;
		#400 //3.4004096e-38 * 7.094076e-33 = 4.7933086e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101011110001011110101011001;
		b = 32'b10111000001001011101000010100001;
		correct = 32'b00100100110000000000001101100110;
		#400 //-3.2920417e-21 * -3.9533366e-05 = 8.3272484e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111100001101010011101111111;
		b = 32'b11000000101110010100000110111100;
		correct = 32'b10111110001110100001001011111011;
		#400 //1.0519866 * -5.789274 = -0.18171303
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000100011000101111111111101;
		b = 32'b10011000101010100000111001011000;
		correct = 32'b00110111010100110101000110001010;
		#400 //-5.5368157e-29 * -4.3958454e-24 = 1.2595565e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100101101001101001001101110;
		b = 32'b11001100101000000010101010001000;
		correct = 32'b00000111100100001000000111101110;
		#400 //-1.8258355e-26 * -83973180.0 = 2.1743078e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100100011100001010010100100;
		b = 32'b11000011110011101011101110001111;
		correct = 32'b11111000001011111111000011000011;
		#400 //5.9017984e+36 * -413.4653 = -1.4273987e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010001010010111101010010110;
		b = 32'b11001111011100011011011001001011;
		correct = 32'b01001010001100110111111100111001;
		#400 //-1.1926014e+16 * -4055255800.0 = 2940878.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001100111000111011001011001;
		b = 32'b00001010111101110100111000000000;
		correct = 32'b11100110001000011111011010101100;
		#400 //-4.553652e-09 * 2.3814575e-32 = -1.9121282e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110100100110100011010001001;
		b = 32'b11011110000111011010110110101000;
		correct = 32'b01011111111011110001110001000100;
		#400 //-9.788138e+37 * -2.8404805e+18 = 3.4459442e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001101111100110101110111111;
		b = 32'b01101100000001111100001000000100;
		correct = 32'b11000101001100111000101000001111;
		#400 //-1.8858371e+30 * 6.564848e+26 = -2872.6287
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000111111100100011111001011110;
		b = 32'b01000000010100000000100010110111;
		correct = 32'b10000111000101010000110001110001;
		#400 //-3.644877e-34 * 3.250532 = -1.121317e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111101001100101110011101100;
		b = 32'b10001010010001110001010111010000;
		correct = 32'b11001100110101011110110001010000;
		#400 //1.0750955e-24 * -9.585604e-33 = -112157310.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110110011000010001101111100011;
		b = 32'b00111000110001001001101001001001;
		correct = 32'b01111101000100101000111100101100;
		#400 //1.1414379e+33 * 9.374746e-05 = 1.2175667e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110011000010110111000010101;
		b = 32'b11010011100011001110101010100101;
		correct = 32'b00000010010011001100010001001111;
		#400 //-1.8210091e-25 * -1210464200000.0 = 1.5043891e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001000110011111101101011010;
		b = 32'b00010110100011111101010110001111;
		correct = 32'b01111010000010010000011111010000;
		#400 //41334186000.0 * 2.323767e-25 = 1.7787578e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110110000110010000011011010;
		b = 32'b10111111101100101100111110011110;
		correct = 32'b01110110100010111010111000111011;
		#400 //-1.9788363e+33 * -1.396961 = 1.4165294e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110001000100111110011001110001;
		b = 32'b01110111011100110011001010111101;
		correct = 32'b00111001000110111010111101111111;
		#400 //7.323661e+29 * 4.9326454e+33 = 0.0001484733
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111010100011011000111111000;
		b = 32'b01011100101110111101010011111001;
		correct = 32'b01100010000011101110011000100001;
		#400 //2.7873272e+38 * 4.229599e+17 = 6.5900505e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101010000000000000001100000;
		b = 32'b11101010001110111001100100011110;
		correct = 32'b00011010100000110000000100100100;
		#400 //-3072.0234 * -5.669805e+25 = 5.418217e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011110110100110010000111000;
		b = 32'b01001001101000011001011001011010;
		correct = 32'b01011001101011001111111100110111;
		#400 //8.0572235e+21 * 1323723.2 = 6086788500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111010101010110011111111001;
		b = 32'b11010111111110110111100100000011;
		correct = 32'b00110110110110010011111110000101;
		#400 //-3580361000.0 * -552994320000000.0 = 6.4744986e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000100010010101001000011011;
		b = 32'b10111101111100000000101000111110;
		correct = 32'b10100010000100100111001101110110;
		#400 //2.3263036e-19 * -0.117207035 = -1.9847814e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001101111010111110111100010001;
		b = 32'b00011000101101111011001111001110;
		correct = 32'b00110100101001000110010011010001;
		#400 //1.4540546e-30 * 4.7485948e-24 = 3.0620734e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101001000100011110110101011;
		b = 32'b01000101111111011010000001011111;
		correct = 32'b10100110101000111100001001011100;
		#400 //-9.222327e-12 * 8116.0464 = -1.1363078e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001111101101000111111010010;
		b = 32'b00010101111011111000111011000100;
		correct = 32'b01110011100000111011111000010000;
		#400 //2019834.2 * 9.6756576e-26 = 2.0875422e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111010001010000011001000011000;
		b = 32'b01011101010010001110011100101111;
		correct = 32'b00011100010101100101001010011111;
		#400 //0.0006416156 * 9.0478695e+17 = 7.0913446e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001010000110010010000000111;
		b = 32'b00011101001110001000110011110100;
		correct = 32'b01010011100001110101100001010111;
		#400 //2.8396714e-09 * 2.4425068e-21 = 1162605400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101011010011101111010010001;
		b = 32'b01011010100010010011101101011110;
		correct = 32'b01010010010110100010001011110000;
		#400 //4.523692e+27 * 1.9313673e+16 = 234222260000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011010000101111110000100010;
		b = 32'b11010111011010000111010110100000;
		correct = 32'b10000011010101101011101100000000;
		#400 //1.6128772e-22 * -255591900000000.0 = -6.3103613e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101000010111001010011001000;
		b = 32'b10110100001111011110100100011011;
		correct = 32'b10110000001111000010011111100101;
		#400 //1.2106737e-16 * -1.76868e-07 = -6.8450695e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001111000001101111111110010;
		b = 32'b11101010100101110010100010101001;
		correct = 32'b00110110101111100110110000001011;
		#400 //-5.1852595e+20 * -9.136991e+25 = 5.675019e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100010110010010011100001000;
		b = 32'b11100010111110111000010111110101;
		correct = 32'b01010000110111010000010001110111;
		#400 //-6.8818363e+31 * -2.3198927e+21 = 29664459000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100010110111100011001010010;
		b = 32'b10100000000000101110000111100000;
		correct = 32'b11101011110101101110111101001100;
		#400 //57612616.0 * -1.1086164e-19 = -5.1968035e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111001110100100011110101110;
		b = 32'b10001010001101100011101101101000;
		correct = 32'b11011100100000101101011111100001;
		#400 //2.5851543e-15 * -8.774154e-33 = -2.9463287e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011111010000100100101011101;
		b = 32'b00111011100010011010010010010000;
		correct = 32'b10001111110110000000001101101000;
		#400 //-8.9473534e-32 * 0.0042005256 = -2.1300556e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101101100001000110100010011;
		b = 32'b10011111100000010101000001000110;
		correct = 32'b01011101101011101100000111110110;
		#400 //-0.08620658 * -5.4766426e-20 = 1.574077e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000011100000001011001011101;
		b = 32'b10110101111101010000000100000111;
		correct = 32'b00011001111110101101110011011001;
		#400 //-4.7348882e-29 * -1.8254221e-06 = 2.5938594e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100010001100011101000011010100;
		b = 32'b00110111000010101111000011100010;
		correct = 32'b11101010101000111101000001000111;
		#400 //-8.2003034e+20 * 8.281526e-06 = -9.9019235e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010101100011000111110110111000;
		b = 32'b11001100011001011001011011101001;
		correct = 32'b10001000100111001010011011111100;
		#400 //5.67439e-26 * -60185508.0 = -9.428166e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111101000011011111010100010;
		b = 32'b00011100000001110010111010100110;
		correct = 32'b01100011000110010010011010110100;
		#400 //1.2636302 * 4.4728045e-22 = 2.8251407e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101100001111001000001110100;
		b = 32'b00100110011101001110001000011101;
		correct = 32'b10011110100011011011011111100110;
		#400 //-1.2748403e-35 * 8.4960946e-16 = -1.5005014e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000000011101001111101111101;
		b = 32'b10000110010011111110010001110011;
		correct = 32'b01110001001011111010000001111011;
		#400 //-3.4003973e-05 * -3.910021e-35 = 8.696622e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000110010000100000000100100;
		b = 32'b11100100100100001011101000110101;
		correct = 32'b11001011101100010001101100011100;
		#400 //4.9579635e+29 * -2.135799e+22 = -23213624.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101100100111010111011011000;
		b = 32'b10011011001001111001001010011111;
		correct = 32'b01101001111000011001110101010001;
		#400 //-4725.8555 * -1.3861292e-22 = 3.4093902e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010011110100011101011000100;
		b = 32'b01000100110111110110100011000111;
		correct = 32'b10011101000011110101110111001100;
		#400 //-3.3912428e-18 * 1787.2743 = -1.8974384e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100010011010101001001101100;
		b = 32'b10111000010001011100100101010110;
		correct = 32'b11100011100001001110000001101111;
		#400 //2.3117198e+17 * -4.715597e-05 = -4.902285e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000110111000100011011000011;
		b = 32'b00110011100111011111111110111111;
		correct = 32'b11111100101100100111001111110001;
		#400 //-5.45378e+29 * 7.357402e-08 = -7.412643e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101111111100001000000110101;
		b = 32'b10101100111001011010010010011000;
		correct = 32'b01111000100011011001110010010001;
		#400 //-1.4997251e+23 * -6.526845e-12 = 2.2977794e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000011011001111011111011100;
		b = 32'b10010101000010101101110000011010;
		correct = 32'b01110010110110100110111110001001;
		#400 //-242655.44 * -2.8042508e-26 = 8.653129e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011010001111010011101111010;
		b = 32'b10110101101101001111100001111110;
		correct = 32'b00111101000011010011011011111101;
		#400 //-4.6485617e-08 * -1.3483366e-06 = 0.03447627
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110000110010010000110101001;
		b = 32'b00111001101101100000001001001100;
		correct = 32'b01011011110101110110001000010100;
		#400 //42092460000000.0 * 0.00034715456 = 1.2124992e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101111010100000111000011001;
		b = 32'b00100101110001110000100101010011;
		correct = 32'b11001111100101101000010100111011;
		#400 //-1.7438462e-06 * 3.4527316e-16 = -5050627600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111001100101110111111101001;
		b = 32'b01000100110001110011110000011111;
		correct = 32'b01100001111001011110101101001110;
		#400 //8.450068e+23 * 1593.8788 = 5.301575e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000111101001011111010111100;
		b = 32'b00001001010001110100001101010001;
		correct = 32'b01110111000111010011011101011010;
		#400 //7.648283 * 2.3985406e-33 = 3.1887237e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011000000011101110011111111;
		b = 32'b01011010010101111011100010110101;
		correct = 32'b01011000000110100001110001011000;
		#400 //1.0288828e+31 * 1.5180052e+16 = 677786100000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010010100000011001000001111101;
		b = 32'b00100011111101000000000101101101;
		correct = 32'b00101110000001111110111011101110;
		#400 //8.176664e-28 * 2.6455137e-17 = 3.090766e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111110000101100101100001010;
		b = 32'b11000000001110101111100011100101;
		correct = 32'b01000111000001010101101010101000;
		#400 //-99734.08 * -2.9214413 = 34138.656
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011101111110100110110100111;
		b = 32'b10111111001010011010100011000001;
		correct = 32'b00000100000100000101010001011010;
		#400 //-1.1243799e-36 * -0.66273123 = 1.6965851e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000010111100011111100011011;
		b = 32'b01111101010110011011001000110110;
		correct = 32'b00100010100000101010110011101110;
		#400 //6.4058194e+19 * 1.8085487e+37 = 3.5419667e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111110000001000010010110001;
		b = 32'b10001110100010011110110110101000;
		correct = 32'b01111111110000001000010010110001;
		#400 //nan * -3.4001962e-30 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100010100001000001100110101;
		b = 32'b01010101100010011011100110111110;
		correct = 32'b01000110010000011100100111001111;
		#400 //2.3476424e+17 * 18928856000000.0 = 12402.452
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011010101001111100010000101;
		b = 32'b00111110101111011111100010010110;
		correct = 32'b10011100000011110111111100110110;
		#400 //-1.761653e-22 * 0.3710372 = -4.7479147e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001101111010110101110011001;
		b = 32'b11011110101000001100010011110001;
		correct = 32'b11011010100101101100111110100110;
		#400 //1.2294081e+35 * -5.7923246e+18 = -2.122478e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101001111100101000110101110;
		b = 32'b00111001010001111110111000010010;
		correct = 32'b00100011011100111011000110011001;
		#400 //2.5188518e-21 * 0.00019066807 = 1.3210664e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001010010010110011100000010;
		b = 32'b11100001101010101001110101000110;
		correct = 32'b10011111000101110001100100011101;
		#400 //12.587648 * -3.934099e+20 = -3.1996267e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111101000110101000100011110;
		b = 32'b10100001001100100101100010000010;
		correct = 32'b11110101111010100110110101100111;
		#400 //359137580000000.0 * -6.0425885e-19 = -5.9434395e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110101110101110111010010011;
		b = 32'b00010110000110110001110011001100;
		correct = 32'b01101000000110100100000111110101;
		#400 //0.36510143 * 1.2529887e-25 = 2.9138445e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111110111010100010011001111;
		b = 32'b01101100110011010110011011001011;
		correct = 32'b10011010100010011110001101010011;
		#400 //-113289.62 * 1.9865218e+27 = -5.7029134e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011101100000000000000111000;
		b = 32'b01000101010001110110001111100100;
		correct = 32'b10000101111000011111100001010111;
		#400 //-6.7793063e-32 * 3190.2432 = -2.1250124e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010011100100111111010110010;
		b = 32'b11100010001011000110111011011100;
		correct = 32'b11010111101101000000001000010100;
		#400 //3.1477638e+35 * -7.9520706e+20 = -395842040000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100010011101010110010010111;
		b = 32'b00101100100010000111100011100001;
		correct = 32'b01000111010000011101100000000111;
		#400 //1.9248033e-07 * 3.8787727e-12 = 49624.027
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100100010100111101001010111;
		b = 32'b00110010111101110101100101011110;
		correct = 32'b11010001000011110101001000110011;
		#400 //-1107.8231 * 2.8795224e-08 = -38472462000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101111110001101010111010010;
		b = 32'b00011010010000111000001110011100;
		correct = 32'b11111011001000101110100010010100;
		#400 //-34199654000000.0 * 4.0431368e-23 = -8.458693e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010110110101001111001000001;
		b = 32'b11000010000001100010111011001010;
		correct = 32'b01011000010100001000101101111100;
		#400 //-3.0767773e+16 * -33.545692 = 917190000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111100001000111000011000001;
		b = 32'b11010111010111001010000011111111;
		correct = 32'b11010111100110011010110001011001;
		#400 //8.1976665e+28 * -242584030000000.0 = -337931000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100111100000010100010010111;
		b = 32'b01010101111111100000011000110100;
		correct = 32'b01011110011100100000011011000111;
		#400 //1.5221857e+32 * 34912824000000.0 = 4.3599614e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101111100111101110100000101;
		b = 32'b10110010000011100010110100001110;
		correct = 32'b11000011010110111000110001100011;
		#400 //1.8169236e-06 * -8.275732e-09 = -219.54839
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001110001111110101111101011;
		b = 32'b00101010010000010001001100000100;
		correct = 32'b00110111000001001000101000011001;
		#400 //1.3547211e-18 * 1.7148441e-13 = 7.8999665e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011101111101110111011001001;
		b = 32'b00111011010010011110100010110001;
		correct = 32'b00011111111100100001010101010011;
		#400 //3.1587175e-22 * 0.003080886 = 1.02526265e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110011101111000101110101010;
		b = 32'b00010000100110010000000011111010;
		correct = 32'b11010101010011110001011101111111;
		#400 //-8.588462e-16 * 6.0349364e-29 = -14231239000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100010000101110011100010111;
		b = 32'b01011011110011111010010010100100;
		correct = 32'b01000111111100000100101011100010;
		#400 //1.438128e+22 * 1.1689269e+17 = 123029.766
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110110011100101000100101011;
		b = 32'b01010111101001011000100010000101;
		correct = 32'b01010110100111111000100101010010;
		#400 //3.192602e+28 * 364011530000000.0 = 87706070000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110110001011101001111100001;
		b = 32'b10111111110101010100000011111110;
		correct = 32'b01010110011011010111101101001100;
		#400 //-108756900000000.0 * -1.6660459 = 65278453000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000000101100010100111000100011;
		b = 32'b10111011111000001010000101011101;
		correct = 32'b10000100010010100001000011100001;
		#400 //1.6282913e-38 * -0.0068551735 = -2.3752736e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100101110010011011001111100;
		b = 32'b01010101000001001111100010110000;
		correct = 32'b10110111001100100100100111001010;
		#400 //-97104860.0 * 9137727000000.0 = -1.0626807e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001000101000010001000011111;
		b = 32'b01111010001010100011110110000010;
		correct = 32'b10010110010111101100000110101000;
		#400 //-39764226000.0 * 2.209845e+35 = -1.7994124e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011011111000001110010111010;
		b = 32'b01111001001100111000011100111100;
		correct = 32'b10101001101100111100000000111010;
		#400 //-4.6506495e+21 * 5.826025e+34 = -7.982543e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010111010111011011110000010;
		b = 32'b11000010010011001111110011000001;
		correct = 32'b01001000000100110011000000111010;
		#400 //-7723969.0 * -51.24683 = 150720.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100011000001101100011110110;
		b = 32'b01001101101011011100010111110100;
		correct = 32'b11000110001001011001111011110010;
		#400 //-3862850700000.0 * 364428930.0 = -10599.736
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000011000110000010011100010001;
		b = 32'b10010000100111101000010000001001;
		correct = 32'b10110001111101011011100100111111;
		#400 //4.471363e-37 * -6.2523444e-29 = -7.1514985e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100111000100011111001101011;
		b = 32'b01011000000000001110101110101010;
		correct = 32'b00110100011000001010000011011001;
		#400 //118616920.0 * 566998600000000.0 = 2.0920142e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011010111010111010101100111;
		b = 32'b10110000001010111110001011110001;
		correct = 32'b10101010101001001110101001001101;
		#400 //1.8318626e-22 * -6.253194e-10 = -2.929483e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111101001011010110000110011;
		b = 32'b11000010001011100011100110000011;
		correct = 32'b10111100111100110110111100011001;
		#400 //1.2943176 * -43.556164 = -0.029716061
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100100011010110010010111001;
		b = 32'b00100000001111000010000101010010;
		correct = 32'b10101011110000000110011100001110;
		#400 //-2.178511e-31 * 1.5935244e-19 = -1.3671024e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011011101010000111010111000;
		b = 32'b10001100011100100001100110101100;
		correct = 32'b11000110100000011001000001000001;
		#400 //3.0930604e-27 * -1.8650727e-31 = -16584.127
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110001111000101010100100000001;
		b = 32'b01111000111000110101000111001100;
		correct = 32'b00111000011111110100000111101001;
		#400 //2.2447336e+30 * 3.68847e+34 = 6.085812e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000001101001011110111111000;
		b = 32'b11011110011111101111001000110010;
		correct = 32'b10000001001101010111110100111111;
		#400 //1.5309448e-19 * -4.5927002e+18 = -3.333431e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011101100111011010110000111;
		b = 32'b10100101000100111100100010000100;
		correct = 32'b10111110000110111010011011101011;
		#400 //1.9484099e-17 * -1.2818155e-16 = -0.15200393
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111001010101111010100110000;
		b = 32'b01110011000101101111111101101001;
		correct = 32'b00110011100100001110101110001000;
		#400 //8.073252e+23 * 1.196327e+31 = 6.7483654e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110000001101101110100111001;
		b = 32'b00001000000001001100100111000011;
		correct = 32'b11000101100000100000000001001100;
		#400 //-1.662329e-30 * 3.9959475e-34 = -4160.037
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000111100110011001011001001;
		b = 32'b00101001001101111011111110100001;
		correct = 32'b11000111001010010110100110111010;
		#400 //-1.7695011e-09 * 4.0800374e-14 = -43369.727
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000101000110001000000010101;
		b = 32'b10100001110111101000111010111010;
		correct = 32'b11111110001110111001000010111011;
		#400 //9.399932e+19 * -1.5081085e-18 = -6.232928e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000110010000110011101010111;
		b = 32'b01011011000100101001001110111000;
		correct = 32'b00111101001011110000000100110101;
		#400 //1762769300000000.0 * 4.1257765e+16 = 0.04272576
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111011101111000110110011111;
		b = 32'b00010111110100010001110100011100;
		correct = 32'b00110111000101111000011101110011;
		#400 //1.22053155e-29 * 1.3513657e-24 = 9.031838e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100001000000111000110001011;
		b = 32'b00110100111101111010101000000010;
		correct = 32'b00111110101001011101100000000000;
		#400 //1.4942468e-07 * 4.6131032e-07 = 0.32391357
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011000111101010111011001101;
		b = 32'b00000010101011000100101001010100;
		correct = 32'b11010111111010111100011111110100;
		#400 //-1.3125935e-22 * 2.531579e-37 = -518488050000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000001011101100000010011001;
		b = 32'b10101001010001100101010010110110;
		correct = 32'b00100110011000011001000011000001;
		#400 //-3.446382e-29 * -4.4038307e-14 = 7.8258735e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100010101111111001100101101;
		b = 32'b11011001000110101100010111011000;
		correct = 32'b11010010101100101001100000110110;
		#400 //1.0442697e+27 * -2722792400000000.0 = -383528930000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011000010110011100110100111;
		b = 32'b10110110110100001011101001111000;
		correct = 32'b10100011101010101100000110010010;
		#400 //1.1516439e-22 * -6.220591e-06 = -1.8513417e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001101110011000100000001000;
		b = 32'b00001100100001111001111101011000;
		correct = 32'b00111100101011110001101010011000;
		#400 //4.4665053e-33 * 2.0895945e-31 = 0.021374986
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000101000000101111110000011;
		b = 32'b01011000101101100101011010100010;
		correct = 32'b01000111011000010010100100111100;
		#400 //9.244879e+19 * 1603865600000000.0 = 57641.234
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101111101111001011101010001;
		b = 32'b11101110100011100010111100011011;
		correct = 32'b10110110110111101110010001010001;
		#400 //1.4615198e+23 * -2.200191e+28 = -6.642695e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111001110010010001011001010;
		b = 32'b01011010101011110000000111111001;
		correct = 32'b10111100000001110110100001100000;
		#400 //-203559070000000.0 * 2.4630145e+16 = -0.008264631
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001000000001110101001010100111;
		b = 32'b00111010110001101001100101000010;
		correct = 32'b10001100101011100110111101111011;
		#400 //-4.072224e-34 * 0.0015151876 = -2.687604e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010101001001101011100001001;
		b = 32'b00011100010111011111010001011010;
		correct = 32'b10110101101111100001111111101101;
		#400 //-1.0402865e-27 * 7.3438583e-22 = -1.4165395e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000011000010110111011001011;
		b = 32'b10010011011011000010011010000100;
		correct = 32'b11000100011101000110000110101000;
		#400 //2.9136505e-24 * -2.9806377e-27 = -977.5259
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110101111100101111111010101;
		b = 32'b00010011010110100101111111011111;
		correct = 32'b01011010110111110010110011101100;
		#400 //8.657223e-11 * 2.7562736e-27 = 3.1409156e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000011000011000110000010000;
		b = 32'b01001011001010001110110001110000;
		correct = 32'b10000100101010101110011111100111;
		#400 //-4.4481326e-29 * 11070576.0 = -4.0179777e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111111101011101010010111010;
		b = 32'b00111000010010000001001100010100;
		correct = 32'b01101111000111010100010111110001;
		#400 //2.3218078e+24 * 4.7701484e-05 = 4.86737e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111100111110011101111000010;
		b = 32'b11110001000111011000011000110110;
		correct = 32'b00110110000000010110001110001010;
		#400 //-1.5039172e+24 * -7.8002236e+29 = 1.9280437e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100000100000111100101111011010;
		b = 32'b01000100101010011100110111110100;
		correct = 32'b11011011010001101011001010111110;
		#400 //-7.597539e+19 * 1358.436 = -5.5928575e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101001101110110111011001100;
		b = 32'b00000100000110010000011100001111;
		correct = 32'b11000000100110010110111010110110;
		#400 //-8.624969e-36 * 1.7988305e-36 = -4.7947645
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011100011001101010101001100;
		b = 32'b10111010000011011000001110001000;
		correct = 32'b11010000111111101100010011001111;
		#400 //18459288.0 * -0.0005398323 = -34194487000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011010111110111011010110000;
		b = 32'b11100101001011100010011011001000;
		correct = 32'b00100101101001000011111001111001;
		#400 //-14644912.0 * -5.1400447e+22 = 2.8491798e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101000101100001010111111101001;
		b = 32'b10100111101111001011001000010000;
		correct = 32'b01000000011011111011010101011010;
		#400 //-1.9616214e-14 * -5.237354e-15 = 3.7454438
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101001010111101100110001111;
		b = 32'b01101001111101111010100111100111;
		correct = 32'b00110010101100011010001001100000;
		#400 //7.739429e+17 * 3.7425877e+25 = 2.0679352e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001000010101111111111000100;
		b = 32'b00011010110101110110011011110110;
		correct = 32'b11100101101001010011001001100101;
		#400 //-8.687443 * 8.908826e-23 = -9.751501e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111010010000001111010101011;
		b = 32'b10000111010011000110101111011010;
		correct = 32'b11010111011110101001110011111000;
		#400 //4.2377015e-20 * -1.5378949e-34 = -275552080000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000010100001011100110011000;
		b = 32'b00111101110110011011101010011110;
		correct = 32'b11010001111101010110100111010000;
		#400 //-14007296000.0 * 0.106312975 = -131755280000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111000010000101000110000110;
		b = 32'b01010101101101111101010011000111;
		correct = 32'b01010000101111011101010110101011;
		#400 //6.437457e+23 * 25265562000000.0 = 25479174000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110001010111011010011111100;
		b = 32'b00011011000000001100100110100001;
		correct = 32'b11100010101010101010100000101001;
		#400 //-0.16768259 * 1.0653062e-22 = -1.5740319e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101111100111011011000111001;
		b = 32'b01010000111001001001110000010100;
		correct = 32'b10001100100010000111010010101110;
		#400 //-6.450998e-21 * 30683472000.0 = -2.1024342e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001101110001001100011010101;
		b = 32'b10101000100111110111101001011101;
		correct = 32'b10111000100101000010100100110111;
		#400 //1.2508779e-18 * -1.7705613e-14 = -7.064867e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101101110110010000111000100;
		b = 32'b10001011010100000001100000110111;
		correct = 32'b11101001111001100011011000100100;
		#400 //1.3942413e-06 * -4.007756e-32 = -3.4788576e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011100111001011101111010101;
		b = 32'b10011010010100010001111100000000;
		correct = 32'b00110000101111111101111001110000;
		#400 //-6.037163e-32 * -4.324523e-23 = 1.39603e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101000011101110000101100111;
		b = 32'b10010100111100111110010000001000;
		correct = 32'b01001111100101011111100101111011;
		#400 //-1.2392906e-16 * -2.4626672e-26 = 5032310300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011100001011000110011000101;
		b = 32'b11010010010011100000010111100111;
		correct = 32'b10011000101001011111001001000011;
		#400 //9.48929e-13 * -221215570000.0 = -4.2896122e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101100101101100110010100010;
		b = 32'b00000101000111000101000101010110;
		correct = 32'b11101111111101101111011001101110;
		#400 //-1.1235427e-06 * 7.350024e-36 = -1.52862455e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011011100101100111000010010;
		b = 32'b01111010011010100110010001100010;
		correct = 32'b10111000100001001001100000011101;
		#400 //-1.9236991e+31 * 3.0425837e+35 = -6.322584e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000010101101100010100110100101;
		b = 32'b00101001000011110010110100110101;
		correct = 32'b10011001001000101101101010000101;
		#400 //-2.67664e-37 * 3.179159e-14 = -8.419333e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101000101010101101100011101001;
		b = 32'b10110010010100100001011011101100;
		correct = 32'b00110101110100000010111010100111;
		#400 //-1.8967861e-14 * -1.2228821e-08 = 1.5510785e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010100001101011010101100110111;
		b = 32'b11000011011000011000010100111000;
		correct = 32'b10010000010011100011100011000110;
		#400 //9.171931e-27 * -225.52039 = -4.0670073e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100010010101011111100011000;
		b = 32'b00101101110010100111001010010101;
		correct = 32'b10100110000000000011000001100000;
		#400 //-1.023608e-26 * 2.3015626e-11 = -4.447448e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101001100010100010001010001;
		b = 32'b11110101100101101010111111001110;
		correct = 32'b00110111000101101001010000001110;
		#400 //-3.4288398e+27 * -3.8203627e+32 = 8.975168e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011101110100000001010010111;
		b = 32'b01001101111000110101110000101110;
		correct = 32'b11010101010100010111000011111001;
		#400 //-6.862562e+21 * 476808640.0 = -14392697000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010000001100110000111001111;
		b = 32'b01011011100010000110001100010001;
		correct = 32'b00101101111111000011110010011100;
		#400 //2201715.8 * 7.677904e+16 = 2.8675999e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000010010111110111110100110;
		b = 32'b11110010000110000111011110110001;
		correct = 32'b10111101101010110011010110000101;
		#400 //2.524607e+29 * -3.019931e+30 = -0.083598174
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010101001011010010111101000;
		b = 32'b00010010100100101010110100000100;
		correct = 32'b01001111100100001000111001111010;
		#400 //4.4899e-18 * 9.256547e-28 = 4850513000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110100101001001111000100100;
		b = 32'b01011111100010010000001010110000;
		correct = 32'b10011110100010101101100000001001;
		#400 //-0.29026902 * 1.9745294e+19 = -1.4700668e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001100110010100110011010011;
		b = 32'b10100111111110100100100000011101;
		correct = 32'b01110001000111001100110101111000;
		#400 //-5393767600000000.0 * -6.9467124e-15 = 7.764489e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010000100001100101000111110;
		b = 32'b11001011001101010110110010110100;
		correct = 32'b00101110010011000100111001111011;
		#400 //-0.00055233005 * -11889844.0 = 4.6453934e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110101000001110100111010101;
		b = 32'b10111111001010000100111110101101;
		correct = 32'b11100110111101001011111101111011;
		#400 //3.7994604e+23 * -0.65746576 = -5.778948e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011011010001011101101010010;
		b = 32'b01100010111011000000010000011011;
		correct = 32'b01001111111111000111000000000110;
		#400 //1.8438907e+31 * 2.1768637e+21 = 8470400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000100111101110010110101101;
		b = 32'b11010110111011011010001001110011;
		correct = 32'b01011001001010110010110101101100;
		#400 //-3.9341034e+29 * -130640985000000.0 = 3011385200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101101111001111010001101110;
		b = 32'b10001001011001011011110111011000;
		correct = 32'b01100011110100101000110100101110;
		#400 //-2.1481674e-11 * -2.7654136e-33 = 7.7679786e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001111000011110001101100011;
		b = 32'b11101011101000110011100100001011;
		correct = 32'b01001101101100010010010001111001;
		#400 //-1.4660984e+35 * -3.9464857e+26 = 371494700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110010101110001110000000110;
		b = 32'b00010010111100001001110111010011;
		correct = 32'b01010010111001001101110010111010;
		#400 //7.463109e-16 * 1.5185036e-27 = 491477860000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111110100000010011000111111;
		b = 32'b10100000101011010111001111110100;
		correct = 32'b11101110100110011001101010110101;
		#400 //6984335000.0 * -2.9384071e-19 = -2.3769118e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000011010000001111110001111;
		b = 32'b00101100110100100010111011100001;
		correct = 32'b01110011000011010101110010000100;
		#400 //6.690498e+19 * 5.9737636e-12 = 1.1199803e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011101001010001110111011100;
		b = 32'b10101101110000111000100010011111;
		correct = 32'b10111101010110000010110101001000;
		#400 //1.1732243e-12 * -2.2229605e-11 = -0.05277756
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010110010000111011011001010;
		b = 32'b11001111011101110010110000000010;
		correct = 32'b01011010110011111001111110110110;
		#400 //-1.21173065e+26 * -4146856400.0 = 2.9220462e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010011101000001010001100001;
		b = 32'b01100110101010100101011001010001;
		correct = 32'b01000011001101110110100111101111;
		#400 //7.3768534e+25 * 4.0219728e+23 = 183.4138
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101010101111101010100101110;
		b = 32'b10101101011100011111001100110011;
		correct = 32'b11001111011001000101110110111001;
		#400 //0.05269354 * -1.3753265e-11 = -3831347500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111111100001000011101010100;
		b = 32'b11100001110101101111100000001110;
		correct = 32'b10110101100011110011100000011000;
		#400 //528928040000000.0 * -4.9568468e+20 = -1.0670656e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100010000100111101010000111;
		b = 32'b00101110010011110010100110011000;
		correct = 32'b11011101011100000101001101110100;
		#400 //-50981404.0 * 4.7103293e-11 = -1.082332e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000001011000001001000011010;
		b = 32'b00111001111011011110100000011001;
		correct = 32'b10010101101110010010100000111000;
		#400 //-3.3934964e-29 * 0.0004537709 = -7.478436e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010110010101010001100111000;
		b = 32'b01011101001001111011000111100011;
		correct = 32'b00101101000110101010101111100100;
		#400 //6640028.0 * 7.5523055e+17 = 8.792054e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011110100001101000011110001;
		b = 32'b00011101111101001010101011111100;
		correct = 32'b11111101010110100111110011011101;
		#400 //-1.1755306e+17 * 6.4763056e-21 = -1.8151252e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110101101101110010000110010;
		b = 32'b11001110110001110110000010000010;
		correct = 32'b00111111011010101101010100011111;
		#400 //-1534204200.0 * -1672495400.0 = 0.91731447
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000111000001111110000010000;
		b = 32'b00001011010100010001011111110111;
		correct = 32'b11001101000010011011101001011010;
		#400 //-5.815716e-24 * 4.0269965e-32 = -144418200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101001011100000110010001100;
		b = 32'b10011011111000010101101110110011;
		correct = 32'b01100000110001011011011011011111;
		#400 //-0.042492434 * -3.7282387e-22 = 1.1397456e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101011011111111011011101001;
		b = 32'b10011101100100000110100000110110;
		correct = 32'b11000111010101001011001101010011;
		#400 //2.0813602e-16 * -3.8224234e-21 = -54451.324
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011111100100110101111101011;
		b = 32'b10100111010111010001110110010010;
		correct = 32'b10111100000011000101010101101110;
		#400 //2.6283398e-17 * -3.0685941e-15 = -0.00856529
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011110111001100100111011000011;
		b = 32'b00000001100000101010010110100000;
		correct = 32'b01011100111000011010010000111010;
		#400 //2.4384772e-20 * 4.799212e-38 = 5.080995e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110111110010011010000110110;
		b = 32'b10110010001110111100001010111011;
		correct = 32'b00111100001010011110001100010110;
		#400 //-1.13324836e-10 * -1.0929109e-08 = 0.010369083
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101101101010010101100101111001;
		b = 32'b11010011001011000111110111101100;
		correct = 32'b10011001111110110101011000011000;
		#400 //1.925281e-11 * -740847000000.0 = -2.5987565e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010110001100101000010000011;
		b = 32'b10001010011000010010010001011111;
		correct = 32'b10110111111000010111111011010101;
		#400 //2.9139697e-37 * -1.08401966e-32 = -2.6881151e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011011100011010101010100000;
		b = 32'b01000011000011011000000111101111;
		correct = 32'b11101111110110101001100100101011;
		#400 //-1.9146793e+31 * 141.50755 = -1.353058e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011110000011011011011100110;
		b = 32'b11000110100010001001111110011101;
		correct = 32'b10001100101101010111110011001010;
		#400 //4.89004e-27 * -17487.807 = -2.796257e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100101001000111110110111110;
		b = 32'b11011010100100101000111100010010;
		correct = 32'b11010001100011111010100101011010;
		#400 //1.5908611e+27 * -2.0626327e+16 = -77127700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100001111111010100110111001;
		b = 32'b11010011010110001000111000110111;
		correct = 32'b01000000011000101001001011001011;
		#400 //-3292745000000.0 * -930098900000.0 = 3.5402095
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000110000100000010011111110;
		b = 32'b10010111101111011001001100111011;
		correct = 32'b00111000100000110000000000110110;
		#400 //-7.65272e-29 * -1.2251005e-24 = 6.246606e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110111110001000000110001010;
		b = 32'b01000110111011110111111010100000;
		correct = 32'b00110111100001001101000011110011;
		#400 //0.4853633 * 30655.312 = 1.5832926e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001110011001001011011101010001;
		b = 32'b01010010000111101111101000111011;
		correct = 32'b00111011101110000010011001010101;
		#400 //959304770.0 * 170700750000.0 = 0.005619804
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000110101111101110110111001;
		b = 32'b10111100010110111101010000010111;
		correct = 32'b01001011111110110110001010111001;
		#400 //-442093.78 * -0.013417265 = 32949618.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011111011000000011100011110011;
		b = 32'b10011100000110101011111001000111;
		correct = 32'b01000010101110010111100010111000;
		#400 //-4.7480952e-20 * -5.1200253e-22 = 92.73578
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110011000111101000001101001;
		b = 32'b11011001011010001100010000011011;
		correct = 32'b01011100011110101000110111000100;
		#400 //-1.1551547e+33 * -4094863400000000.0 = 2.8209847e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100101111010011000000000010;
		b = 32'b00110011110101010001110001111000;
		correct = 32'b11001000011000110100001011111101;
		#400 //-0.023094181 * 9.923764e-08 = -232715.95
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101111101110001101001110000;
		b = 32'b10110000001100010011110110100000;
		correct = 32'b00101101001100100111010000010101;
		#400 //-6.540769e-21 * -6.44798e-10 = 1.0143904e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110000011010101011111001001;
		b = 32'b00001010011111010001111000010101;
		correct = 32'b11100011000011101111001111011000;
		#400 //-3.2137657e-11 * 1.2187165e-32 = -2.6370085e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111000111110010111000010011;
		b = 32'b00111100011000000110111001110001;
		correct = 32'b01010010001101011001000111111110;
		#400 //2670596900.0 * 0.013698206 = 194959600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110011101110011110010011101;
		b = 32'b01000101010011001100101100110111;
		correct = 32'b01010000100110101000011100010100;
		#400 //67959926000000.0 * 3276.701 = 20740350000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010001100110101111110000101;
		b = 32'b01111010010010101101010111110101;
		correct = 32'b10110111011000100110001100111111;
		#400 //-3.5528507e+30 * 2.6329588e+35 = -1.3493757e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011100000011011001011010111;
		b = 32'b00110100110111101111000010001101;
		correct = 32'b11010110000101001110111010010101;
		#400 //-16999854.0 * 4.1525746e-07 = -40938106000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111111000101010000000101011;
		b = 32'b10110000100001111110110100100111;
		correct = 32'b11111110110101010110100100000111;
		#400 //1.4027449e+29 * -9.889946e-10 = -1.4183545e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111001111001010111101110010;
		b = 32'b11000100101010101000110111010010;
		correct = 32'b00111010000011011001101110000101;
		#400 //-0.7370521 * -1364.4319 = 0.00054018974
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110000010001011110011111110;
		b = 32'b10101110100011001000111110110100;
		correct = 32'b11001110111110010000100110000001;
		#400 //0.13353345 * -6.39199e-11 = -2089074800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101100111001001011010100011;
		b = 32'b11100100111010101000110101101000;
		correct = 32'b00110000001010101110100000110000;
		#400 //-21521350000000.0 * -3.461382e+22 = 6.21756e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001010001100101011111011111;
		b = 32'b10001000100011001001001110111101;
		correct = 32'b11011000001101001001100100010011;
		#400 //6.7201306e-19 * -8.460677e-34 = -794278200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111101100100110110101110010;
		b = 32'b10001111001110111110011011110100;
		correct = 32'b11101111111100110001011101110110;
		#400 //1.393965 * -9.264292e-30 = -1.5046644e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100100010100101000001010001;
		b = 32'b10111101110110100000111011000111;
		correct = 32'b10111110001000100110000101100111;
		#400 //0.016884001 * -0.1064735 = -0.15857469
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010110010110000100000011111;
		b = 32'b11111000100011110100010010110001;
		correct = 32'b10111001101101010110010011110010;
		#400 //8.042915e+30 * -2.3246615e+34 = -0.0003459822
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000101110100000100011010011;
		b = 32'b10111011111010111000001001011110;
		correct = 32'b10010100010010100011100001111010;
		#400 //7.337766e-29 * -0.007187172 = -1.0209532e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000010111100111110001101000;
		b = 32'b11111110011000110000110111100001;
		correct = 32'b10000001011110101101100101110000;
		#400 //3.4763432 * -7.5451705e+37 = -4.6073752e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011001000000101011111011111;
		b = 32'b11011100101011100111010010111011;
		correct = 32'b10001101111010110100101001101100;
		#400 //5.6965365e-13 * -3.9283994e+17 = -1.450091e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110001101001011011110011011;
		b = 32'b01010010001110100110101000010110;
		correct = 32'b01101011011110000010110100010111;
		#400 //6.0053593e+37 * 200160940000.0 = 3.0002653e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011011110110100001010001000;
		b = 32'b01101100100100110011000000000001;
		correct = 32'b01000110010110101000000101100001;
		#400 //1.9906859e+31 * 1.4235103e+27 = 13984.345
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000110110010101011000011000;
		b = 32'b11100101100110111110010100000001;
		correct = 32'b10111010101100100111001010100110;
		#400 //1.2528585e+20 * -9.20239e+22 = -0.001361449
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111110010010010001110100110;
		b = 32'b10111110010000011010101000101000;
		correct = 32'b11011001000001001111000010110010;
		#400 //442309900000000.0 * -0.18912566 = -2338709000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100001011001001111111111011;
		b = 32'b11000100100101011001101110010110;
		correct = 32'b11001111000100111011000101011100;
		#400 //2965673600000.0 * -1196.862 = -2477874200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111000010110010000000011010;
		b = 32'b10100011001010110001101100100011;
		correct = 32'b11100011010100000010011011111011;
		#400 //35616.1 * -9.275675e-18 = -3.8397316e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110011010111101011111010011;
		b = 32'b01000011111010000011101110011101;
		correct = 32'b00110010000000011111110101100110;
		#400 //3.5143355e-06 * 464.46573 = 7.566404e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000010101110100100111000010001;
		b = 32'b00101111101100011100011100011001;
		correct = 32'b10010010100001100010001110111101;
		#400 //-2.7375052e-37 * 3.233758e-10 = -8.465399e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000010011011000000010111011;
		b = 32'b01000100001010100111110110100000;
		correct = 32'b00010011100110100100100101000100;
		#400 //2.6560621e-24 * 681.9629 = 3.894731e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110110110111100010110001010;
		b = 32'b00101001000100100001001111110100;
		correct = 32'b00111101010000001001001011011110;
		#400 //1.5249721e-15 * 3.243582e-14 = 0.047015063
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110010010101010101110111000;
		b = 32'b01110110110110110110110011101110;
		correct = 32'b10010110111011000111001111011010;
		#400 //-850062850.0 * 2.225239e+33 = -3.820097e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110111110001101110100111110;
		b = 32'b10100110101010010100100011111110;
		correct = 32'b11000111101111000010101111100010;
		#400 //1.1317035e-10 * -1.1746515e-15 = -96343.766
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100010011110000110110111001101;
		b = 32'b11111011000000011111110011001010;
		correct = 32'b00100110111101001010000101101010;
		#400 //-1.1456761e+21 * -6.749335e+35 = 1.6974652e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100000110000011110111101101;
		b = 32'b10011011100111100110111010010111;
		correct = 32'b11010111111101011111111101110010;
		#400 //1.4178632e-07 * -2.6210374e-22 = -540954960000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100100110110010000000011000;
		b = 32'b10011001100110101011101100010001;
		correct = 32'b01111010100000000101001110010011;
		#400 //-5330067000000.0 * -1.5998782e-23 = 3.3315454e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100110000111010101011001000;
		b = 32'b11100011110110001001011001110011;
		correct = 32'b11000000011001110100010111000100;
		#400 //2.887537e+22 * -7.9906755e+21 = -3.6136332
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001001000011000100000111110;
		b = 32'b01000110100001101011010010110101;
		correct = 32'b01001010000110010111110110101000;
		#400 //43360970000.0 * 17242.354 = 2514794.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110000001010000000010111101;
		b = 32'b11110011101001101110001011111011;
		correct = 32'b10111001110011000000010111101101;
		#400 //1.02906e+28 * -2.6444244e+31 = -0.00038914327
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110101001011111001010010010;
		b = 32'b01101101000100001001011011000001;
		correct = 32'b00001001000100101110100001111100;
		#400 //4.945622e-06 * 2.7967557e+27 = 1.7683424e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101111111101111111111100001101;
		b = 32'b10110110100110001010100101101001;
		correct = 32'b00111000110011111110111100000111;
		#400 //-4.5110263e-10 * -4.549675e-06 = 9.9150515e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100101000011100111001000010;
		b = 32'b11100011111011101000100001111001;
		correct = 32'b01011000001011011010011101110101;
		#400 //-6.7211456e+36 * -8.800318e+21 = 763738940000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100000111111100111100100101;
		b = 32'b01101100101101101001100000100001;
		correct = 32'b11001110111000000000111000010001;
		#400 //-3.3191064e+36 * 1.7659433e+27 = -1879509100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010111111010010001111000111;
		b = 32'b01110001110100100110001011110011;
		correct = 32'b00010000100110100000001011100001;
		#400 //126.56988 * 2.0835672e+30 = 6.0746725e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011111010110010011111011011;
		b = 32'b01111111011000111100110110111101;
		correct = 32'b00011100000001000010000110001010;
		#400 //1.3238088e+17 * 3.02803e+38 = 4.3718485e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011100110011101010001100100100;
		b = 32'b11011010000011000101111001010000;
		correct = 32'b10000010001111000110110111111110;
		#400 //1.3674107e-21 * -9877549000000000.0 = -1.3843625e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111000011001101100001100001;
		b = 32'b01011111000000101111100110010111;
		correct = 32'b01001111100010011010010101100101;
		#400 //4.3589487e+28 * 9.43774e+18 = 4618636000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011110101101000000011100000;
		b = 32'b10100000001011100110010000110101;
		correct = 32'b11001011000111010111000100000010;
		#400 //1.5241385e-12 * -1.4771529e-19 = -10318082.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010100000010001000110110100;
		b = 32'b00111001000010001000100011011010;
		correct = 32'b00111000111100100000000010100001;
		#400 //1.5025627e-08 * 0.00013020952 = 0.000115395764
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110101000100011100110111001;
		b = 32'b11100001011001110100000011001110;
		correct = 32'b11001100101100111001010111100111;
		#400 //2.5103177e+28 * -2.6661672e+20 = -94154550.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010111011110101001111001100;
		b = 32'b11010011011111110001001000110100;
		correct = 32'b11100110111100000011001011101011;
		#400 //6.2132928e+35 * -1095522060000.0 = -5.671536e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110010011110101000000010111;
		b = 32'b01110000011111011110110000001011;
		correct = 32'b11000101010100010000001001100111;
		#400 //-1.05120104e+33 * 3.1434026e+29 = -3344.1501
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111010100101101010111110101;
		b = 32'b01100001101010101110101101111100;
		correct = 32'b11000101000111011110010010000000;
		#400 //-9.956438e+23 * 3.9411437e+20 = -2526.2812
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010101000111010110101010101101;
		b = 32'b00010111111110101101100111100000;
		correct = 32'b10111100101000001010010111010111;
		#400 //-3.179005e-26 * 1.6210871e-24 = -0.019610329
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110100101101110000010011110;
		b = 32'b01011111100101110101100100100011;
		correct = 32'b10000110011111110011010000100101;
		#400 //-1.0469223e-15 * 2.1811573e+19 = -4.799848e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110001011000010110000101011;
		b = 32'b01011000100011000101011100011111;
		correct = 32'b10110101000111010000100001111101;
		#400 //-722143940.0 * 1234446500000000.0 = -5.849941e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100001100011110101110111011;
		b = 32'b00011011110100011110101011010001;
		correct = 32'b01000111110110001111101010111101;
		#400 //3.858043e-17 * 3.4727896e-22 = 111093.48
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101111101000010011010010110111;
		b = 32'b00001001110011101001011000111011;
		correct = 32'b01100101010001111100001110110110;
		#400 //2.9323186e-10 * 4.9733972e-33 = 5.8960072e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100010111100110010100111111;
		b = 32'b11001011110110000101001000001010;
		correct = 32'b11011000000000111001100000111101;
		#400 //1.6409891e+22 * -28353556.0 = -578759500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110101101101000010000110011001;
		b = 32'b01110000111101001110011010011010;
		correct = 32'b11000100001111000100101110000110;
		#400 //-4.5668695e+32 * 6.0634498e+29 = -753.18005
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110100001111010010010110010001;
		b = 32'b01010111110001011010111100101101;
		correct = 32'b10011011111101001111000110100110;
		#400 //-1.7615663e-07 * 434712330000000.0 = -4.0522576e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010010111011110111001100010;
		b = 32'b10100001111101001110101111011011;
		correct = 32'b11001111111001111111100001001110;
		#400 //1.2918095e-08 * -1.6596514e-18 = -7783619600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111000100100111000000110000;
		b = 32'b11000001110111110111011111010110;
		correct = 32'b10001100101001111100000110011110;
		#400 //7.219962e-30 * -27.933514 = -2.5846953e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001110110100011000100010101;
		b = 32'b10101110010100111100000001001001;
		correct = 32'b01111011000000111110010010101100;
		#400 //-3.2972202e+25 * -4.814663e-11 = 6.848289e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110001101011000101101101100;
		b = 32'b01110101101001101100000001111110;
		correct = 32'b10001000000010110101101011100000;
		#400 //-0.17728966 * 4.2276635e+32 = -4.1935614e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000110000101001101100101110;
		b = 32'b01110000101100011011100110011000;
		correct = 32'b10011111100011000010100001110111;
		#400 //-26119598000.0 * 4.4002573e+29 = -5.935925e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111011100111001011001101110;
		b = 32'b00010011101100100001011100011000;
		correct = 32'b11111011001011110001001101001101;
		#400 //-4086722000.0 * 4.495629e-27 = -9.090434e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001111100010111101101101111;
		b = 32'b00100100010110101100001001001101;
		correct = 32'b11001101000011010100101110110111;
		#400 //-7.028056e-09 * 4.7435794e-17 = -148159340.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000100011101100110010101001110;
		b = 32'b01000000101110111011001000010101;
		correct = 32'b00000011001010000000011111100100;
		#400 //2.8963678e-36 * 5.8654885 = 4.937982e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000001010101100101011010111;
		b = 32'b11011000011010001110101101111100;
		correct = 32'b00110111001110111011011101011011;
		#400 //-11461680000.0 * -1024392400000000.0 = 1.1188759e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101100011101101111100001010010;
		b = 32'b10010101110110001111101110101001;
		correct = 32'b01010110000100011011000010000110;
		#400 //-3.5096548e-12 * -8.7638755e-26 = 40046837000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100100010101001110010110110011;
		b = 32'b10000000000000100001101011101100;
		correct = 32'b01100110010010100100001100010000;
		#400 //-4.6164735e-17 * -1.93329e-40 = 2.3878878e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101010111100010111010010101;
		b = 32'b00100011010010010000010000011111;
		correct = 32'b00100001100011010111101001001001;
		#400 //1.04469456e-35 * 1.08971045e-17 = 9.5869e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101111100010110011101001111;
		b = 32'b10000001110010101111101011101110;
		correct = 32'b11000011100110000011101011011011;
		#400 //2.270148e-35 * -7.456315e-38 = -304.4598
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000001101000000100000000110;
		b = 32'b01110010110011010010001001101010;
		correct = 32'b10110100111000001010110000011100;
		#400 //-3.400696e+24 * 8.126212e+30 = -4.1848477e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100001000100000000011011111;
		b = 32'b10100111101000100011001001100101;
		correct = 32'b11011011111111111011000111010110;
		#400 //648.0136 * -4.501867e-15 = -1.439433e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000001000011000001111111110;
		b = 32'b11011001001010111110101011110100;
		correct = 32'b00110110011100001000001010100001;
		#400 //-10839128000.0 * -3024409700000000.0 = 3.5838823e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110010101111000010001111000;
		b = 32'b00101011010011101100010011010110;
		correct = 32'b10100010100001010110101001110001;
		#400 //-2.6564577e-30 * 7.3459067e-13 = -3.616242e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110101111011000101101100000;
		b = 32'b01001101100111101100110001000110;
		correct = 32'b11011000100110001100100010001100;
		#400 //-4.4754914e+23 * 333023420.0 = -1343896900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000011101001001000111001000101;
		b = 32'b10011101001000010111111001111001;
		correct = 32'b01100110000000100110110100111101;
		#400 //-329.11148 * -2.1373557e-21 = 1.5398068e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111001000101110000110101011101;
		b = 32'b10001010000101111001011101010011;
		correct = 32'b01101110011111110001011100000101;
		#400 //-0.0001440546 * -7.2988465e-33 = 1.9736627e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000111001000011011001100101;
		b = 32'b11001001011110110010011111110101;
		correct = 32'b10001110111010001001110100101000;
		#400 //5.8991543e-24 * -1028735.3 = -5.734375e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101000101010110011001001000;
		b = 32'b11001101110111110100000010100111;
		correct = 32'b00111110101010110101000001100001;
		#400 //-156656770.0 * -468194530.0 = 0.33459762
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001110010011111000110010001;
		b = 32'b10110010110111000000000001011010;
		correct = 32'b01001110011010101111110011001011;
		#400 //-25.242952 * -2.561153e-08 = 985608900.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000011010011101000011111100;
		b = 32'b11111101001110001010001001010011;
		correct = 32'b00011010101000100001100010100100;
		#400 //-1028335160000000.0 * -1.5338799e+37 = 6.704144e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110011000000000110100011101;
		b = 32'b10110000001111011100011010111100;
		correct = 32'b11110101100101110001111000100001;
		#400 //2.64513e+23 * -6.904022e-10 = -3.8312886e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111010111100000010011011110;
		b = 32'b11001001010110001111010000101100;
		correct = 32'b01011101100000101111110100001001;
		#400 //-1.04845514e+24 * -888642.75 = 1.1798388e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011100010110001111000100010;
		b = 32'b01101000111000111010011111001011;
		correct = 32'b01001010000111000111000001010010;
		#400 //2.204408e+31 * 8.6005794e+24 = 2563092.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101000111110011000000100001100;
		b = 32'b00100010010110110101010100010100;
		correct = 32'b11000110000100011001101110100000;
		#400 //-2.7700518e-14 * 2.9725074e-18 = -9318.906
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000100001011100011100010001;
		b = 32'b00010111101011101011010001000011;
		correct = 32'b11011000010001000000011101101000;
		#400 //-9.733602e-10 * 1.1289991e-24 = -862144350000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011110001001100000110100011101;
		b = 32'b11000011110001101010111111001100;
		correct = 32'b10011001110101011111001101010010;
		#400 //8.7906786e-21 * -397.3734 = -2.212196e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101001000011100100101001011;
		b = 32'b01001011011101001111000001110110;
		correct = 32'b00111001001010010001011110010010;
		#400 //2588.5808 * 16052342.0 = 0.00016125877
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001001010111111001101000000;
		b = 32'b01010100111001010001011000110011;
		correct = 32'b00101011110000000010011010101010;
		#400 //10.746887 * 7871359600000.0 = 1.3653152e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111001100101101100000101010;
		b = 32'b11010010000010100110001011000011;
		correct = 32'b01010100101001010110110000010110;
		#400 //-8.4456876e+23 * -148590610000.0 = 5683864000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000101011011100000010010010;
		b = 32'b11110011100011111111001110001001;
		correct = 32'b10010100100110100111111110101001;
		#400 //355844.56 * -2.2809995e+31 = -1.5600379e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011011010110000101010111101;
		b = 32'b11010001010000111101001011111001;
		correct = 32'b11011001100110011010001001111001;
		#400 //2.8414828e+26 * -52566135000.0 = -5405539000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110100101111101100001001111;
		b = 32'b00001110100101110111100110110100;
		correct = 32'b01011111100000000100111111110010;
		#400 //6.905109e-11 * 3.734157e-30 = 1.849175e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010011000010110110110100000;
		b = 32'b01101100100000010101110001010000;
		correct = 32'b10101101010111110000111010100101;
		#400 //-1.5863101e+16 * 1.2510989e+27 = -1.2679334e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100001010110001000111011011;
		b = 32'b00101010100100110000110100000010;
		correct = 32'b11101001000101001110100001000000;
		#400 //-2938956000000.0 * 2.6121472e-13 = -1.1251112e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101000010100110010010101101;
		b = 32'b11000001010101101101011101101000;
		correct = 32'b10011011001001001110011111111010;
		#400 //1.8316196e-21 * -13.427589 = -1.3640718e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101111100110110110010010011;
		b = 32'b00111101111011001111101110111111;
		correct = 32'b10111111100000110111101010010010;
		#400 //-0.11885943 * 0.11571454 = -1.027178
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111010011101010111001001000;
		b = 32'b01001101011010011111010100000101;
		correct = 32'b10110001011000100010011101011101;
		#400 //-0.8073468 * 245321810.0 = -3.2909704e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100011100100001100101000110;
		b = 32'b10110101000010111010110111100010;
		correct = 32'b01001110110111011101101100010001;
		#400 //-968.3949 * -5.203457e-07 = 1861060700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001110111110011010001101000;
		b = 32'b10110000000000101101101000101010;
		correct = 32'b01010001010110100101011011101001;
		#400 //-27.900589 * -4.7603754e-10 = 58610060000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101011000110101101110011110;
		b = 32'b00110000010110000110000010001000;
		correct = 32'b11101100100001100111111011101101;
		#400 //-1.02392886e+18 * 7.871752e-10 = -1.3007636e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111101010010101100001010111;
		b = 32'b00000010111100101001001111011110;
		correct = 32'b01111100001100101011011100100001;
		#400 //1.3230084 * 3.5643576e-37 = 3.7117725e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001100110101100011100101000;
		b = 32'b01111110000100111001101101010010;
		correct = 32'b00001011000001100011011111111011;
		#400 //1267941.0 * 4.9050746e+37 = 2.5849576e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001110010100001010011000111;
		b = 32'b11010101001100000000101000001011;
		correct = 32'b10111100000100101110111101110100;
		#400 //108491500000.0 * -12097324000000.0 = -0.008968223
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010011111011000100001100001;
		b = 32'b00111011101010001101110111010100;
		correct = 32'b10100110010000000010110100110100;
		#400 //-3.4360092e-18 * 0.005153397 = -6.6674643e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000011100001110000110011100;
		b = 32'b10100011111110001011010001010100;
		correct = 32'b11100011111101111111001010001000;
		#400 //246662.44 * -2.6964586e-17 = -9.147644e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000110010111111001011000100;
		b = 32'b00100000001111001000110110111000;
		correct = 32'b01110000000010100111001101100011;
		#400 //27373478000.0 * 1.597111e-19 = 1.713937e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001011100100111110001000001;
		b = 32'b00011001011011001111111100010100;
		correct = 32'b01001111100000101111011011101101;
		#400 //5.3842567e-14 * 1.2252427e-23 = 4394441000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110011100110011010100011001;
		b = 32'b10000011000001101101100101011101;
		correct = 32'b11111010111001101101101011010001;
		#400 //0.23750724 * -3.962858e-37 = -5.993332e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110001101110011001101011111;
		b = 32'b01110001000010101111110010000111;
		correct = 32'b00001100101010001011100000100000;
		#400 //0.1789069 * 6.882275e+29 = 2.5995315e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010001100101111000101110101;
		b = 32'b01101011110010001000010101101110;
		correct = 32'b11000101111001000111001110110010;
		#400 //-3.544335e+30 * 4.8483054e+26 = -7310.462
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101000001100001000011110101010;
		b = 32'b00010000001100100110111001111010;
		correct = 32'b11010111011111010100010110001111;
		#400 //-9.79938e-15 * 3.5189418e-29 = -278475200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010100111001101010001000110001;
		b = 32'b01010011011011011110100100100101;
		correct = 32'b00000000111110000010101101100110;
		#400 //2.3288038e-26 * 1021818770000.0 = 2.2790771e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011001001100111011001011000;
		b = 32'b10010111100000001110010100110000;
		correct = 32'b11000011001001010100111001011100;
		#400 //1.3769437e-22 * -8.329661e-25 = -165.30609
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100101111100010111010110100;
		b = 32'b10110101010100110100010001101100;
		correct = 32'b11101110111001100111001101100101;
		#400 //2.8065974e+22 * -7.870319e-07 = -3.5660528e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100101000011010010111101100;
		b = 32'b01001100110100100000111111011100;
		correct = 32'b01011111010001001111111110101000;
		#400 //1.5633648e+27 * 110132960.0 = 1.4195249e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001110100001111100110011011;
		b = 32'b10100010110000010111000011010101;
		correct = 32'b10101110100010100100011101110000;
		#400 //3.2970445e-28 * -5.243222e-18 = -6.288203e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000010100110100100101101000;
		b = 32'b11011000101000011101000111011010;
		correct = 32'b00100111001001110010000011101011;
		#400 //-3.3013554 * -1423381400000000.0 = 2.319375e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111011111000110001100000100;
		b = 32'b01000001110001101101000100110011;
		correct = 32'b00001101001000100111110100001111;
		#400 //1.2443629e-29 * 24.852148 = 5.007064e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010001111001100000001111110;
		b = 32'b11111011010110010010101000010110;
		correct = 32'b10110110010111101000000110101011;
		#400 //3.738617e+30 * -1.127582e+36 = -3.3156055e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000011011011101000111101101;
		b = 32'b01010010000100110001111110110110;
		correct = 32'b11011101110011101110100000110011;
		#400 //-2.9440693e+29 * 157973050000.0 = -1.8636528e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101101100011000110111101001;
		b = 32'b11111111000001100011011011111010;
		correct = 32'b10001110001010010101010100110000;
		#400 //372358430.0 * -1.78402e+38 = -2.0871875e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100000001101010101010010110;
		b = 32'b10101110100111101001010011110011;
		correct = 32'b01011100110110010110010010011110;
		#400 //-35301976.0 * -7.211467e-11 = 4.895256e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010011111111000001100010000;
		b = 32'b00011001000101100101000110100100;
		correct = 32'b11000000110110011001001100000101;
		#400 //-5.2838635e-23 * 7.7713054e-24 = -6.7991967
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111100000001100010110011101;
		b = 32'b10111011110111101101010101010001;
		correct = 32'b01100011000100111111000001000000;
		#400 //-1.855799e+19 * -0.0068003316 = 2.7289832e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001101000011100001011101111;
		b = 32'b00110001000011110000011100111111;
		correct = 32'b01011000000100001100001111001011;
		#400 //1325149.9 * 2.0813358e-09 = 636682400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100001100000011001110010100;
		b = 32'b11001010000001111010010011110111;
		correct = 32'b00000001101001100100010101111101;
		#400 //-1.3574068e-31 * -2222397.8 = 6.107848e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110001100110110111101010011;
		b = 32'b00111011000111110100101110100010;
		correct = 32'b00011010100100000010111011001100;
		#400 //1.4494633e-25 * 0.0024306555 = 5.963261e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100001011011000011011000100;
		b = 32'b11010010010011110011011000101010;
		correct = 32'b01000001010101100110001000110100;
		#400 //-2981161300000.0 * -222491740000.0 = 13.398975
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011100111011100110111111011;
		b = 32'b10101111111000111101111001100111;
		correct = 32'b11111011001100010100100101000011;
		#400 //3.8154814e+26 * -4.1449086e-10 = -9.205225e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101010101100010010011011000;
		b = 32'b00000010111001000111100101111101;
		correct = 32'b11011001111011111111000101100000;
		#400 //-2.8341712e-21 * 3.357132e-37 = -8442239000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111101011101011101101011000;
		b = 32'b01010000101010111010001110010000;
		correct = 32'b01000110100000100100111001111001;
		#400 //384239320000000.0 * 23036985000.0 = 16679.236
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010100111111100001101110100100;
		b = 32'b10100110011011000100111001010101;
		correct = 32'b10101110000010011010010010001111;
		#400 //2.5658348e-26 * -8.198511e-16 = -3.129635e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000001101111110101000100010;
		b = 32'b01001001111111111000001001111101;
		correct = 32'b11100101101110000100010001111010;
		#400 //-2.2767522e+29 * 2093135.6 = -1.08772325e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000001001111100000001110011;
		b = 32'b01010111011101111001101011001101;
		correct = 32'b00111000001011010111000010000111;
		#400 //11257630000.0 * 272244240000000.0 = 4.1351213e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100110011100111000001011010;
		b = 32'b11010000101110110000001101000001;
		correct = 32'b00001011100011010100101111010000;
		#400 //-1.3660979e-21 * -25100421000.0 = 5.4425294e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011110100101110110111000101;
		b = 32'b11101001000010010011010010110010;
		correct = 32'b11001010010001001100011011001001;
		#400 //3.3423e+31 * -1.036698e+25 = -3223986.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100110111010101011111111010;
		b = 32'b00001000011000100001110111010000;
		correct = 32'b01011011111110101001100010110000;
		#400 //9.599251e-17 * 6.8044446e-34 = 1.4107325e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101000101110101110110111010;
		b = 32'b11001010110001010011111001101000;
		correct = 32'b10010001110001000111010010111110;
		#400 //2.003314e-21 * -6463284.0 = -3.0995295e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010110011011110000101011110;
		b = 32'b10011101100010010101001011000100;
		correct = 32'b01101100101111111110011100001001;
		#400 //-6746287.0 * -3.6349176e-21 = 1.8559669e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000000110000111000001100010;
		b = 32'b11111000001011000001100110000000;
		correct = 32'b00110111011000101100000100101111;
		#400 //-1.8871034e+29 * -1.3962379e+34 = 1.3515629e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110011100011101000000100100;
		b = 32'b00101011000010001101011100010110;
		correct = 32'b10110010111000100011000011111111;
		#400 //-1.2801476e-20 * 4.86154e-13 = -2.6332144e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110000101100100111110001110;
		b = 32'b00011000010011111111101001010001;
		correct = 32'b01010101001110010000010010000010;
		#400 //3.417671e-11 * 2.68805e-24 = 12714313000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011100111100011011011111101001;
		b = 32'b01011000101011010010000110100011;
		correct = 32'b00000011101100101011010100111100;
		#400 //1.5995582e-21 * 1522879800000000.0 = 1.0503509e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001001011110111011100000000;
		b = 32'b01010110111010101111010100100001;
		correct = 32'b00110001101111110010110111100010;
		#400 //718704.0 * 129169270000000.0 = 5.564048e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100010101111111001111100101;
		b = 32'b10010100101010001010100100010100;
		correct = 32'b00111111001000111110010000011111;
		#400 //-1.0902826e-26 * -1.7030354e-26 = 0.6401996
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100010010100010111001000110;
		b = 32'b01001001110101110000100000110110;
		correct = 32'b01100001111100001011001101000011;
		#400 //9.7768614e+26 * 1761542.8 = 5.5501697e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101001010110000110110010011;
		b = 32'b01110110000010010000000110000111;
		correct = 32'b00001110100111111100111100011011;
		#400 //2736.8484 * 6.947028e+32 = 3.939596e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001100111101111010100010101;
		b = 32'b11010111100000011010111111110100;
		correct = 32'b01000001100111001110001110100011;
		#400 //-5592814600000000.0 * -285185430000000.0 = 19.61115
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000011001010010111100010000000;
		b = 32'b00101001010101001010011110011010;
		correct = 32'b11011001010011000000001110001011;
		#400 //-169.4707 * 4.7218827e-14 = -3589049400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010110111101111100011001110;
		b = 32'b10111111110101110011101011100000;
		correct = 32'b00010010100001001001101010101110;
		#400 //-1.4071505e-27 * -1.6814842 = 8.368503e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110111011100110110010000010;
		b = 32'b00011011100100001100110100101000;
		correct = 32'b01100010110100101100001001101000;
		#400 //0.4656716 * 2.395538e-22 = 1.9439124e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001111111011101101110011110;
		b = 32'b00010011111010110010111110101001;
		correct = 32'b11101101100010100010100101111101;
		#400 //-31.732235 * 5.9369337e-27 = -5.344886e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011101111100110101010100011;
		b = 32'b01110110110100010111001001111101;
		correct = 32'b01000100011010001011110101001110;
		#400 //1.9773985e+36 * 2.1240472e+33 = 930.9579
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000001111110001101011101111;
		b = 32'b01111011000111000100011111011001;
		correct = 32'b10001100100111001000010111001110;
		#400 //-195691.73 * 8.1145555e+35 = -2.4116136e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010011011110001100111000101;
		b = 32'b01010100001111000010011010001001;
		correct = 32'b00000101101000101010100101100101;
		#400 //4.9444858e-23 * 3232401500000.0 = 1.5296633e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110101101011110011001010001;
		b = 32'b01101101011001010010001100100101;
		correct = 32'b00110000110010110011100101111011;
		#400 //6.5536264e+18 * 4.4321596e+27 = 1.4786531e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000010001110001111110111010;
		b = 32'b10001101101001011101001000111111;
		correct = 32'b01110010000110011011010011110011;
		#400 //-3.1113114 * -1.0219525e-30 = 3.0444775e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101110010101010111011100011;
		b = 32'b00101001001010000111001000000111;
		correct = 32'b10111100000110100000010001010100;
		#400 //-3.5159922e-16 * 3.7402397e-14 = -0.009400446
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011000011010011001011001011;
		b = 32'b00110000110100011111011000000010;
		correct = 32'b11011001101011000010100011011011;
		#400 //-9253579.0 * 1.5276671e-09 = -6057327000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001000100011010111100000101;
		b = 32'b11100011110110101101111101110111;
		correct = 32'b00101100101010100110010101010010;
		#400 //-39106662000.0 * -8.074985e+21 = 4.8429394e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100100100000000011001100000;
		b = 32'b01000010100101100111001100010101;
		correct = 32'b10011001011101010001000101101100;
		#400 //-9.530769e-22 * 75.22477 = -1.26697214e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010011001111111110111000100;
		b = 32'b01011010001001100111001110100111;
		correct = 32'b00111111101100100110011000111010;
		#400 //1.6324934e+16 * 1.1713002e+16 = 1.3937447
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111111001101110001011110011;
		b = 32'b00110110011110101100110100011111;
		correct = 32'b11101000111010111010110000100111;
		#400 //-3.3274254e+19 * 3.73723e-06 = -8.903454e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011001111001111001111100010111;
		b = 32'b00100011111110100010101100100101;
		correct = 32'b10110101011011010000010101000100;
		#400 //-2.3949096e-23 * 2.7123327e-17 = -8.829704e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111100011110010000000000010;
		b = 32'b10101011100111110110101011110101;
		correct = 32'b11010011011001011101011000011100;
		#400 //1.1181643 * -1.1327316e-12 = -987139700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101111010000000101001111000;
		b = 32'b00110010001101001111101010101100;
		correct = 32'b11000011001001000001110100110101;
		#400 //-1.7288394e-06 * 1.0534375e-08 = -164.11409
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010000010110011100011110000;
		b = 32'b00010110101100011000101010111110;
		correct = 32'b00110010110010001011111100011110;
		#400 //6.703315e-33 * 2.868345e-25 = 2.3369974e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101000011010110010111010110;
		b = 32'b00110000010011111001010111101000;
		correct = 32'b01010100001011100110000000100000;
		#400 //2262.3647 * 7.551919e-10 = 2995748000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001110110000011110111111001;
		b = 32'b00110101000110101100110001100001;
		correct = 32'b01100100001100101100111010000101;
		#400 //7608342000000000.0 * 5.766688e-07 = 1.3193607e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011001011000001101110111110;
		b = 32'b01011110100111110111100111101011;
		correct = 32'b01011100000010100010001110001110;
		#400 //8.936377e+35 * 5.745737e+18 = 1.5553056e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010010100101110000110111110000;
		b = 32'b11010110011111011110010101011000;
		correct = 32'b00111011100110000100111001101001;
		#400 //-324386950000.0 * -69790366000000.0 = 0.004648019
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110010101011001010010000010;
		b = 32'b00111011011010110011001001011000;
		correct = 32'b10111010011010000111100010110001;
		#400 //-3.1825916e-06 * 0.0035888162 = -0.0008868082
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111110111010010101000110001;
		b = 32'b10111100101000111110110110100101;
		correct = 32'b01011010101011001011000100100011;
		#400 //-486346560000000.0 * -0.020010779 = 2.430423e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010001001011111100110000101;
		b = 32'b11001111111000111110011100000010;
		correct = 32'b10111001101110100110111111111000;
		#400 //2719329.2 * -7647134700.0 = -0.00035560108
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011001001000111000101000010;
		b = 32'b01001110110001011001000110000101;
		correct = 32'b11101011110101010001001110101100;
		#400 //-8.538338e+35 * 1657324200.0 = -5.151882e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010011000010000001010001001;
		b = 32'b11011001110011111101010010011011;
		correct = 32'b01011000000010101001010010100000;
		#400 //-4.4567803e+30 * -7312385300000000.0 = 609483800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111000000100110010100100001001;
		b = 32'b10010110000001000011101111001011;
		correct = 32'b11100001100011100111001011100111;
		#400 //3.5085748e-05 * -1.0681742e-25 = -3.2846466e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010001010110101111000001010;
		b = 32'b10100100011010111011010000101001;
		correct = 32'b10110101001110100001111110100111;
		#400 //3.5437935e-23 * -5.1110104e-17 = -6.933646e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011010001011011010101101000;
		b = 32'b01011000100100100011000101010110;
		correct = 32'b00010010001011010001101011100111;
		#400 //7.024021e-13 * 1285924800000000.0 = 5.4622334e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001110011010100000111110011;
		b = 32'b10111011110101001101001111001111;
		correct = 32'b11001101011101101110010100001010;
		#400 //1681470.4 * -0.006494976 = -258887840.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011111000011111111000100100;
		b = 32'b01111000110110011000111000110111;
		correct = 32'b10011010100001001111011011001110;
		#400 //-1941262800000.0 * 3.5300402e+34 = -5.4992655e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101010100001111000100100111;
		b = 32'b00010011001111001100101011000010;
		correct = 32'b01010001100011011010100101011101;
		#400 //1.812283e-16 * 2.3828903e-27 = 76053980000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110001101110101001101010100;
		b = 32'b10110111011100110001001000000011;
		correct = 32'b01011110010000010001001110111111;
		#400 //-50392130000000.0 * -1.4488122e-05 = 3.4781684e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100001001011100110000110000;
		b = 32'b10100101100001101001110101011000;
		correct = 32'b01110110000111011010011010010110;
		#400 //-1.8667151e+17 * -2.3351915e-16 = 7.9938415e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110110100111111111110101000111;
		b = 32'b00111000001110110011111100111101;
		correct = 32'b01111101110110101011101111100011;
		#400 //1.6224849e+33 * 4.464317e-05 = 3.6343408e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100111010100010111000111111;
		b = 32'b01011111010110100100001001111010;
		correct = 32'b10101101000010010101011001000100;
		#400 //-122778104.0 * 1.5727267e+19 = -7.806703e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011111111100000110101010100100;
		b = 32'b00110101100110111111000000110010;
		correct = 32'b10101001110001010101011111001101;
		#400 //-1.01820376e-19 * 1.1618306e-06 = -8.7637884e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100010010110000000011011001100;
		b = 32'b00101110011110101101001100110000;
		correct = 32'b11110011010111000111101111001111;
		#400 //-9.962466e+20 * 5.703099e-11 = -1.7468513e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110000011101010000000011100;
		b = 32'b11001111010110110001001010011101;
		correct = 32'b01100110001001101010101010101000;
		#400 //-7.231968e+32 * -3675430100.0 = 1.9676522e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111011101000110101000011010;
		b = 32'b00110101000011011101000110101101;
		correct = 32'b11100001110111001001100100101111;
		#400 //-268736540000000.0 * 5.283171e-07 = -5.086652e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001100011111101111011110011;
		b = 32'b11001111011000000100111100100100;
		correct = 32'b00100001101001000011001010000000;
		#400 //-4.187194e-09 * -3763283000.0 = 1.112644e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000101010010010001001000011;
		b = 32'b11111110101010000010000110010000;
		correct = 32'b10000001100000001100001101101110;
		#400 //5.2854323 * -1.1174228e+38 = -4.73002e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000110101001000101101000011;
		b = 32'b00111110110100111010000111101011;
		correct = 32'b01010001100000001000110100100010;
		#400 //28527172000.0 * 0.4133447 = 69015450000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001010001011001001110010110;
		b = 32'b00001111010111111001100111100101;
		correct = 32'b10111001011000100011010001011010;
		#400 //-2.3782407e-33 * 1.1024388e-29 = -0.00021572542
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111110110011101110111100011;
		b = 32'b00010110011100001101000011100101;
		correct = 32'b00110000111001111001101010001111;
		#400 //3.2780944e-34 * 1.9452961e-25 = 1.685139e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010010000000101101100100101;
		b = 32'b10110011010111001110010000100010;
		correct = 32'b11110110010111101110110111110001;
		#400 //5.8136044e+25 * -5.1430227e-08 = -1.13038665e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001101000001111010101100110;
		b = 32'b10111010001101010000001000010001;
		correct = 32'b00001110111000111010010011011100;
		#400 //-3.874937e-33 * -0.000690491 = 5.6118574e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101111110010111010111111100;
		b = 32'b00110100010011100100101100000001;
		correct = 32'b01111001000110101100100011100000;
		#400 //9.65055e+27 * 1.9212531e-07 = 5.0230497e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101101110110000110010100010;
		b = 32'b10011111001110101101010011011000;
		correct = 32'b11111110000000000010011000111001;
		#400 //1.6847907e+18 * -3.9563092e-20 = -4.258491e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001110011011001101001110010;
		b = 32'b11111110010101001001100000111001;
		correct = 32'b00010010111101111001010011001110;
		#400 //-110382430000.0 * -7.064668e+37 = 1.5624575e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000000000110011011010110000100;
		b = 32'b00111010000001011000001110000001;
		correct = 32'b00000100110001010010110111000011;
		#400 //2.361003e-39 * 0.0005093143 = 4.6356503e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101000000011100111010110001;
		b = 32'b10001000010111011101001110111101;
		correct = 32'b00111100000101011100110111110010;
		#400 //-6.103514e-36 * -6.6753666e-34 = 0.0091433395
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101101011111101101011101010;
		b = 32'b01111101110000100010001100111100;
		correct = 32'b10100111011001111110010001001001;
		#400 //-1.0380655e+23 * 3.2256647e+37 = -3.2181443e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100000110010101101110011001;
		b = 32'b11101111101011010011000010001110;
		correct = 32'b00011011111000101010111110000001;
		#400 //-40201828.0 * -1.0719921e+29 = 3.750198e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010100000110110101111101000;
		b = 32'b00101001011101010011010110000010;
		correct = 32'b00011000100010010011010001111100;
		#400 //1.9310655e-37 * 5.444734e-14 = 3.5466666e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010111101110000101011001110;
		b = 32'b00111010011011001100100100101010;
		correct = 32'b01010000000001011000101101011010;
		#400 //8095079.0 * 0.00090326613 = 8962009000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100110011011111100111001101;
		b = 32'b10101011010100001110101011001101;
		correct = 32'b11001000111111000110010101001101;
		#400 //3.836598e-07 * -7.4222296e-13 = -516906.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111001000001010100111111010;
		b = 32'b01110100111110010010101101110010;
		correct = 32'b10111001101001010001000101110001;
		#400 //-4.972309e+28 * 1.57930065e+32 = -0.00031484247
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010011010001011101000111010011;
		b = 32'b01111000100011000110101111000100;
		correct = 32'b00011010001101000101001001001011;
		#400 //849628800000.0 * 2.2784603e+34 = 3.7289603e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101010100010010010011101000;
		b = 32'b10111001010100110001010010000011;
		correct = 32'b00001011011111011010011011101101;
		#400 //-9.8339114e-36 * -0.0002013017 = 4.885161e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110111101101011110011101000;
		b = 32'b01001110000110001001010010010101;
		correct = 32'b11011000010011101111110100101010;
		#400 //-5.8259343e+23 * 639968600.0 = -910346900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000011101010010011001011111;
		b = 32'b00011100011101111011011010010001;
		correct = 32'b11010011011111010101100111011010;
		#400 //-8.918501e-10 * 8.1961406e-22 = -1088134200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100111100001011010110000101;
		b = 32'b10110101101001011101011111110000;
		correct = 32'b11000110101110011100100000111010;
		#400 //0.02938343 * -1.2356304e-06 = -23780.113
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001000101101001001011001011;
		b = 32'b01011010100011100100010000111001;
		correct = 32'b11001110000001110111100101010001;
		#400 //-1.1377005e+25 * 2.002223e+16 = -568218700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001110010110101011110001011;
		b = 32'b11000010011111000101100010100000;
		correct = 32'b01101110110011100100100101000110;
		#400 //-2.0138013e+30 * -63.086548 = 3.1921247e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110001011000000101001010010000;
		b = 32'b01110001111011001111110111110110;
		correct = 32'b00111110111100100101000001110111;
		#400 //1.1107913e+30 * 2.3470554e+30 = 0.47327015
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101100101101001010001110000010;
		b = 32'b10000011010010001100100001110001;
		correct = 32'b11101000111001100101000011011110;
		#400 //5.1340607e-12 * -5.9004813e-37 = -8.701088e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100110110111101010110011010;
		b = 32'b11001111000011011010001011100101;
		correct = 32'b11010101010001101010101101011110;
		#400 //3.2441829e+22 * -2376263000.0 = -13652457000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110010110001010111001000100;
		b = 32'b00110010100000101010000011100111;
		correct = 32'b11011011010101000101001000010110;
		#400 //-908824800.0 * 1.5207162e-08 = -5.976295e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011101001100110101000110011;
		b = 32'b01100110110010010001011001011011;
		correct = 32'b00111100010100111101101111110100;
		#400 //6.139624e+21 * 4.7480402e+23 = 0.012930859
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100111010001001000010100000;
		b = 32'b11000010111010100101010010000111;
		correct = 32'b11110001011111100001001001001111;
		#400 //1.4740554e+32 * -117.16509 = -1.2581012e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101000010110101011111011001;
		b = 32'b11001111110011110110010011111100;
		correct = 32'b00011100101011000000000000000000;
		#400 //-7.920741e-12 * -6959003600.0 = 1.1382005e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100001010100010100110101000011;
		b = 32'b00011000111111000000101011000110;
		correct = 32'b11000111110101001001011010101011;
		#400 //-7.091421e-19 * 6.515135e-24 = -108845.336
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101000011101010000100110111110;
		b = 32'b10100111110101111001000011010001;
		correct = 32'b01000000000100011000000000010011;
		#400 //-1.36023446e-14 * -5.9831498e-15 = 2.273442
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000011010110101000111110011;
		b = 32'b01000010111100100010010001011001;
		correct = 32'b01011100111110001100100110100111;
		#400 //6.7826405e+19 * 121.07099 = 5.602201e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101010100100111111111110110;
		b = 32'b00000110100111101001100001010000;
		correct = 32'b01101110001010011110010001001011;
		#400 //7.8417304e-07 * 5.96568e-35 = 1.3144739e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101101011110101100011001001;
		b = 32'b10010011001110100000101011001110;
		correct = 32'b01011001111100010100100001100110;
		#400 //-1.9934625e-11 * -2.3481828e-27 = 8489384000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010101001000100101101111100;
		b = 32'b10110111010111000100010100100000;
		correct = 32'b01100010101111101111000111110011;
		#400 //-2.3122446e+16 * -1.3129116e-05 = 1.7611578e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110110011011100100000101000;
		b = 32'b00001001011010010000010111011110;
		correct = 32'b11100100111000100001001010100111;
		#400 //-9.3578756e-11 * 2.8049114e-33 = -3.3362466e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101010101111010000110011110;
		b = 32'b11011101100011000011010110101010;
		correct = 32'b10110111010001001101101010011000;
		#400 //14818071000000.0 * -1.262896e+18 = -1.1733406e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011000110100010010110101110;
		b = 32'b10000011100010001110111100010001;
		correct = 32'b01110111000100000001011100011110;
		#400 //-0.0023520994 * -8.0482485e-37 = 2.9224985e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111010011101101010011101100110;
		b = 32'b10101001000100100001101001100010;
		correct = 32'b11010000110110000001011110001100;
		#400 //0.00094090996 * -3.2441396e-14 = -29003375000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101111111001101110100001110;
		b = 32'b01101100101110111000100111100101;
		correct = 32'b00001000101011001001010111111110;
		#400 //1.8839798e-06 * 1.8137625e+27 = 1.0387136e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111000001101111000001010011;
		b = 32'b11001010001100011001010011101011;
		correct = 32'b10011100010000101000011011000000;
		#400 //1.8726516e-15 * -2909498.8 = -6.4363376e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010001010001111101111001001;
		b = 32'b11110011000001010000001000011001;
		correct = 32'b11000110101000101001111011101010;
		#400 //2.1935317e+35 * -1.0537995e+31 = -20815.457
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100000100010000101100011011101;
		b = 32'b01100001010101011010000011001011;
		correct = 32'b10111110101000110110010000001011;
		#400 //-7.8598765e+19 * 2.4629643e+20 = -0.31912264
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001010100101111101111001100;
		b = 32'b01001110101100111010111011011000;
		correct = 32'b01011010000101100100110000100111;
		#400 //1.5941469e+25 * 1507290100.0 = 1.0576244e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010100110000110001100000000;
		b = 32'b11000111111011100000011001101000;
		correct = 32'b01101010001000111110010100000000;
		#400 //-6.03666e+30 * -121868.81 = 4.9534083e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000110111011110111110001011010;
		b = 32'b00010000110010000111010100011110;
		correct = 32'b10110101100110001110101111001100;
		#400 //-9.0084526e-35 * 7.906654e-29 = -1.1393508e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001101010101100000100000011;
		b = 32'b11110111001111110010101100001001;
		correct = 32'b00111001111001001010100110100101;
		#400 //-1.6910652e+30 * -3.8773498e+33 = 0.00043613944
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101010100000011000111101111;
		b = 32'b10010010010011000001101111110010;
		correct = 32'b11001010100000101000111111110101;
		#400 //2.7554386e-21 * -6.4405495e-28 = -4278266.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011011101100111000110111100;
		b = 32'b10010010000010010011011111010110;
		correct = 32'b01101000111001011110001101110110;
		#400 //-0.0037604412 * -4.32984e-28 = 8.6849427e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100000100111101101001101010;
		b = 32'b10101011010100010001001001001100;
		correct = 32'b01111000001101010000101001100001;
		#400 //-1.0909639e+22 * -7.427711e-13 = 1.4687754e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001010100100000000100011010;
		b = 32'b00101101100000010111011000000101;
		correct = 32'b11010011010011111010001001100011;
		#400 //-13.125269 * 1.4718013e-11 = -891782600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011011010111101100000010000;
		b = 32'b11000011011101110010111101111101;
		correct = 32'b11010111011101000100000100001010;
		#400 //6.6384183e+16 * -247.1855 = -268560180000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101010111011000100010001101;
		b = 32'b00010111111111000101011110111111;
		correct = 32'b01011100111000001011111001111111;
		#400 //8.2527623e-07 * 1.6307269e-24 = 5.0607878e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110111111110101100001000101;
		b = 32'b01100100100111001110110001100101;
		correct = 32'b00000001110100000100011111100011;
		#400 //1.7718105e-15 * 2.3157809e+22 = 7.6510285e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001101110010011001100110001100;
		b = 32'b11000000001111011101100010010110;
		correct = 32'b10001101000001111110110010111100;
		#400 //1.2424546e-30 * -2.9663444 = -4.1885045e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111001110111011010011110100;
		b = 32'b11111000000111010010001010011000;
		correct = 32'b00110110100110001110011100111101;
		#400 //-5.8092456e+28 * -1.2748316e+34 = 4.5568727e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000101110000110010000000101;
		b = 32'b11110010100100101111010010011100;
		correct = 32'b00001101101000001001101101000100;
		#400 //-5.7622094 * -5.8215073e+30 = 9.89814e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101001000001000100010000010001;
		b = 32'b10100000010010110100001101111101;
		correct = 32'b01001000001001101001010100000000;
		#400 //-2.9368926e-14 * -1.7217099e-19 = 170580.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000011001110111001110110010;
		b = 32'b01000111000110000010010000101101;
		correct = 32'b11100000110000101011100111010010;
		#400 //-4.3720034e+24 * 38948.176 = -1.1225182e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010100010111100110011110000;
		b = 32'b00100111011111010110000100010101;
		correct = 32'b01001010100011010011111100011101;
		#400 //1.6274925e-08 * 3.5163431e-15 = 4628366.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111001011010000000001001110100;
		b = 32'b01010100000001000100010011001001;
		correct = 32'b00100100111000001000010110011111;
		#400 //0.00022126158 * 2272358800000.0 = 9.737088e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001110000011110111110111101;
		b = 32'b11101111100001010011100000100100;
		correct = 32'b00100001101110100101011010100000;
		#400 //-104118850000.0 * -8.245875e+28 = 1.262678e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110001000001101000010000001;
		b = 32'b00111011101010010100011100001111;
		correct = 32'b01000001111100110011001110000000;
		#400 //0.15704538 * 0.0051659415 = 30.400146
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101100001000011001100010110;
		b = 32'b10100100010000010000101100111101;
		correct = 32'b01000000101011110101000000011010;
		#400 //-2.2932967e-16 * -4.1859723e-17 = 5.478528
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110110001101010101001101001;
		b = 32'b01111010001111001000101001101010;
		correct = 32'b10000100000001101101111110110100;
		#400 //-0.38801888 * 2.447398e+35 = -1.5854344e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011100111110111011000000110;
		b = 32'b00000110011110110010111001101000;
		correct = 32'b11110100101000101000010100101010;
		#400 //-0.0048663644 * 4.7241947e-35 = -1.030094e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010011110110010010110111001;
		b = 32'b01101001110100000100100010000011;
		correct = 32'b00100000000110100101011110010000;
		#400 //4114798.2 * 3.1474875e+25 = 1.307328e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110101100010011111000010010101;
		b = 32'b11001011011101000000110010010101;
		correct = 32'b01101001100100001011000111001110;
		#400 //-3.4971887e+32 * -15994005.0 = 2.1865622e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100011111010100010111001100;
		b = 32'b10010110001011000010100011010011;
		correct = 32'b11111101101111000100111010110000;
		#400 //4351191000000.0 * -1.3906931e-25 = -3.128793e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100101001111110101001011111;
		b = 32'b10111000001110000011110110010100;
		correct = 32'b01111011111010010101000100001011;
		#400 //-1.064291e+32 * -4.3926368e-05 = 2.4228978e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000010111111100000111101001;
		b = 32'b00000011011010000101011000011011;
		correct = 32'b11011100011101101000110000011111;
		#400 //-1.8952994e-19 * 6.8277517e-37 = -2.7758764e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101000110101001011111000010111;
		b = 32'b11001010111000110011100110100110;
		correct = 32'b10011101011011111010111011101111;
		#400 //2.3619166e-14 * -7445715.0 = -3.1721825e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000101000111000000111111001;
		b = 32'b11110001000101010100100100010100;
		correct = 32'b00110111000011000011000111000100;
		#400 //-6.1771465e+24 * -7.392258e+29 = 8.356237e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011111010011010001111001001;
		b = 32'b01100011011010110110000110111110;
		correct = 32'b00100111111111100001101011111011;
		#400 //30623634.0 * 4.342028e+21 = 7.0528414e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110111111001111000001110000;
		b = 32'b11100010111100101110000000101011;
		correct = 32'b10011011100001010100110110111110;
		#400 //0.4940219 * -2.2401325e+21 = -2.2053244e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101010000111000001101000010;
		b = 32'b00100110001000011011011010000100;
		correct = 32'b01001110100110101100000011011111;
		#400 //7.2834166e-07 * 5.610545e-16 = 1298165600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001010101001110011001010110;
		b = 32'b11000101001011001010111001010101;
		correct = 32'b00101011100111011100111111101101;
		#400 //-3.098099e-09 * -2762.8958 = 1.1213232e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101010000110110011011100000;
		b = 32'b00000010000101000110111110100101;
		correct = 32'b01000010101010000111111111101011;
		#400 //9.187751e-36 * 1.0905363e-37 = 84.24984
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000110001101101110011110001110;
		b = 32'b00000110001111001101011100100100;
		correct = 32'b10111111011101111111001111111100;
		#400 //-3.4400515e-35 * 3.551693e-35 = -0.96856666
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111010111110110111100010110;
		b = 32'b01001011010111110111001011111100;
		correct = 32'b00000011011111111111101110001001;
		#400 //1.1016143e-29 * 14643964.0 = 7.5226513e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011100101010001011010110000;
		b = 32'b01110110101111111111001101000001;
		correct = 32'b11000100010001101101011000011110;
		#400 //-1.5482248e+36 * 1.9466064e+33 = -795.3456
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110001111000010011101110110;
		b = 32'b00000010001001101100010011111001;
		correct = 32'b11110011100100000110100111010001;
		#400 //-2.8037152e-06 * 1.2252282e-37 = -2.2883208e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110101000111011000110100000;
		b = 32'b00111101101101110100111110111000;
		correct = 32'b00001000011001001001101001111110;
		#400 //6.157478e-35 * 0.08950752 = 6.879286e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110100010011110011001110101;
		b = 32'b10110101001111011110001111000101;
		correct = 32'b00100000101110011110100100001010;
		#400 //-2.2278983e-25 * -7.0739435e-07 = 3.1494431e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101011010100010111110000110;
		b = 32'b00100101100111001110001100110011;
		correct = 32'b10110111001111110001000010111010;
		#400 //-3.0994211e-21 * 2.7215642e-16 = -1.1388382e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001011000111001110001011101;
		b = 32'b11001000010001000111010110000010;
		correct = 32'b10000000100101000100101111100111;
		#400 //2.7397653e-33 * -201174.03 = -1.3618882e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010001111111010111010100101;
		b = 32'b00000010011100010010110000110110;
		correct = 32'b11101111010010110111011110000010;
		#400 //-1.1157373e-08 * 1.7718572e-37 = -6.2969933e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001101101011111000111101010100;
		b = 32'b11001100011010011101101001011010;
		correct = 32'b00000000110000000010111110110001;
		#400 //-1.0819713e-30 * -61303144.0 = 1.7649524e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010101001100100100110000001;
		b = 32'b01001010000111110100001101000001;
		correct = 32'b00101000000001011010010101000011;
		#400 //1.935837e-08 * 2609360.2 = 7.4188185e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011000110110011101101111111;
		b = 32'b11101010111111101110100010011000;
		correct = 32'b10110111100110111110010110100110;
		#400 //2.8635325e+21 * -1.5408278e+26 = -1.8584378e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101101100001001101011101001;
		b = 32'b10010001010100110110011101101010;
		correct = 32'b11110011110101011101110000111011;
		#400 //5651.364 * -1.6676832e-28 = -3.3887513e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110110010001100111100000100;
		b = 32'b11001111001111000110111111011000;
		correct = 32'b00101111000010000110011101011111;
		#400 //-0.3922044 * -3161446400.0 = 1.2405853e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111001010011000010001111001110;
		b = 32'b00111111000111100001110001010110;
		correct = 32'b00111001101001010100001101101011;
		#400 //0.00019468294 * 0.6176199 = 0.00031521483
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110010100011001011010001111;
		b = 32'b00110110100001100000100000111111;
		correct = 32'b01001111010010000010011111001100;
		#400 //13413.64 * 3.994471e-06 = 3358051300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010100011010110010001100100;
		b = 32'b11011100000100101110001010010001;
		correct = 32'b11001101111101100110110100111100;
		#400 //8.546631e+25 * -1.6537784e+17 = -516794240.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111000000110011001011110010;
		b = 32'b10101000111101000111000111011000;
		correct = 32'b10100101100010010110011010101000;
		#400 //6.46861e-30 * -2.7138814e-14 = -2.3835274e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111100001000111110000010111;
		b = 32'b11001101111000101111100111111111;
		correct = 32'b10000001000101010110110011101111;
		#400 //1.3064003e-29 * -476004320.0 = -2.7445134e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001000101110011110010111101;
		b = 32'b11111110010110110001111010010110;
		correct = 32'b00111010001100001011000100111111;
		#400 //-4.9079297e+34 * -7.2814936e+37 = 0.0006740279
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001110111111111100110010101;
		b = 32'b01101101011000100110000011001101;
		correct = 32'b10101011111111010100100001000111;
		#400 //-7880417300000000.0 * 4.3787898e+27 = -1.7996792e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101100010001110101000100010;
		b = 32'b10000111010101100101111011010100;
		correct = 32'b01111101101000111000000010101110;
		#400 //-4381.2666 * -1.6127438e-34 = 2.7166538e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110110101101111001110011101;
		b = 32'b10100011111010011110010110010100;
		correct = 32'b11100010011010110100001110110111;
		#400 //27513.807 * -2.535914e-17 = -1.08496606e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111111011100000010011011100;
		b = 32'b01001001001001010111010110101000;
		correct = 32'b11001110001110000010000111010100;
		#400 //-523409280000000.0 * 677722.5 = -772306200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111010100111001010101110111;
		b = 32'b00100011001110011110011001001001;
		correct = 32'b01111011100100011010111101001101;
		#400 //1.5246223e+19 * 1.0077635e-17 = 1.5128771e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000011011011100001101010110;
		b = 32'b10101110111001000110010011011100;
		correct = 32'b11110001000001010100000000110001;
		#400 //6.853053e+19 * -1.0386156e-10 = -6.5982574e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000001001001011110001010001;
		b = 32'b11010101010011011010110001000111;
		correct = 32'b00101010010011010000101110100110;
		#400 //-2.573994 * -14133738000000.0 = 1.8211699e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010100010001000111011111000;
		b = 32'b01010100111101110101000001111100;
		correct = 32'b00110101000011010101101010111000;
		#400 //4474748.0 * 8497658000000.0 = 5.2658606e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000101010001100110100100111;
		b = 32'b01001000110010011101011100111001;
		correct = 32'b10100111010101100001100001100111;
		#400 //-1.2281917e-09 * 413369.78 = -2.9711694e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110010001110110100111010111;
		b = 32'b10101000111000011000010001011111;
		correct = 32'b11111100111000100101111000110011;
		#400 //2.3542583e+23 * -2.5037425e-14 = -9.4029574e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011101110000111100011100000;
		b = 32'b10101011000101000100110001000101;
		correct = 32'b10100000000111110011100100010101;
		#400 //7.1056094e-32 * -5.268601e-13 = -1.3486711e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011101010110101110100101101;
		b = 32'b01110001001000010010000110111011;
		correct = 32'b00001010000010000010000011010110;
		#400 //0.0052296133 * 7.978858e+29 = 6.5543376e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110111101101101000001100000110;
		b = 32'b00111000110111101111001110110001;
		correct = 32'b11111110010100011001000011000011;
		#400 //-7.4035586e+33 * 0.00010631176 = -6.9640074e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011000010010110111100001111;
		b = 32'b00111001100001100100111101011001;
		correct = 32'b10110001000000101111101000100100;
		#400 //-4.88263e-13 * 0.0002561759 = -1.9059678e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010000001100101010110101111;
		b = 32'b00011000100101111000001110001010;
		correct = 32'b11001000111000101111100101010001;
		#400 //-1.8205747e-18 * 3.9165406e-24 = -464842.53
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001110001101110100010011010;
		b = 32'b00010111100011001110111011101010;
		correct = 32'b10101001101101001010011110101111;
		#400 //-7.306748e-38 * 9.107598e-25 = -8.022694e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111111101010001111001001101;
		b = 32'b01011000000000011100001011001011;
		correct = 32'b10110111011100011100101011000001;
		#400 //-8224807400.0 * 570694500000000.0 = -1.4411927e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111101101101101110001100100;
		b = 32'b00110100101001100000101001100001;
		correct = 32'b11101010100011001111011101111101;
		#400 //-2.6353033e+19 * 3.092746e-07 = -8.520917e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110001110001000000110111111;
		b = 32'b00000111011110111100101101001111;
		correct = 32'b01011110001110111001011010110110;
		#400 //6.4013663e-16 * 1.8942888e-34 = 3.3792979e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101111001011011010101010100;
		b = 32'b10101001110010111000001101111110;
		correct = 32'b11001011100100000111100110100011;
		#400 //1.7114603e-06 * -9.037821e-14 = -18936646.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011110110001000010111001001;
		b = 32'b01110010001111100011111111101011;
		correct = 32'b10000001000100011010110100101010;
		#400 //-1.0082619e-07 * 3.768283e+30 = -2.6756533e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010010101001101110010010001;
		b = 32'b11000010010001101001110100100001;
		correct = 32'b11011111100010010010111010100111;
		#400 //9.816508e+20 * -49.653446 = -1.9770044e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101100100110010011000111101;
		b = 32'b00011110011100101111000110110011;
		correct = 32'b00111110100110110000111010100101;
		#400 //3.8950113e-21 * 1.28613556e-20 = 0.3028461
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011001100000000110101110101;
		b = 32'b10011111010011100100101111111110;
		correct = 32'b01011011010110100111100000001110;
		#400 //-0.002686349 * -4.3685056e-20 = 6.1493546e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111110101010110000111101010;
		b = 32'b01001111100011000000110100111001;
		correct = 32'b11000111110000110000010101000110;
		#400 //-469233030000000.0 * 4699353600.0 = -99850.55
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011011101110011001111101011;
		b = 32'b10100010110110011001111110010000;
		correct = 32'b11101000000100010110010111011010;
		#400 //16200683.0 * -5.898691e-18 = -2.746488e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101111111111110110100011000110;
		b = 32'b10100001010010110001010110000010;
		correct = 32'b01001110001000001111101011001000;
		#400 //-4.6458676e-10 * -6.880754e-19 = 675197440.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001101111100001001100111011;
		b = 32'b01011001100010100001101101011000;
		correct = 32'b11000111101100000010101001001011;
		#400 //-4.382834e+20 * 4859201400000000.0 = -90196.586
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000100100000001001000011100;
		b = 32'b11001011101100001001001000001001;
		correct = 32'b11010100010100001110000101100011;
		#400 //8.305113e+19 * -23143442.0 = -3588538200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100110101011100010001110000;
		b = 32'b01111001001001000101111011111100;
		correct = 32'b01000011001001100111011101011000;
		#400 //8.8795477e+36 * 5.334145e+34 = 166.46619
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001100101100111110101101100;
		b = 32'b11011111010001010100010001110111;
		correct = 32'b00101001110000110100101110011111;
		#400 //-1232813.5 * -1.4214617e+19 = 8.672858e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010100100111010110111010000010;
		b = 32'b11000111011000101010001010111111;
		correct = 32'b10001100101100011101010001010111;
		#400 //1.5896536e-26 * -58018.746 = -2.7398965e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110100011011010100100001111011;
		b = 32'b10011010011011010000011111001000;
		correct = 32'b01011001100000000010001011110000;
		#400 //-2.2098713e-07 * -4.9016737e-23 = 4508401400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100001001011111011111100110;
		b = 32'b00111001000110101101110111100001;
		correct = 32'b11000010100010010010110011111010;
		#400 //-0.010129904 * 0.00014769241 = -68.587845
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101100111001100111111000100100;
		b = 32'b00101000001101011101001110100101;
		correct = 32'b11000100001000100100001001011110;
		#400 //-6.5509976e-12 * 1.00934115e-14 = -649.037
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110100111110110111011111101;
		b = 32'b00001111011101110101000101000000;
		correct = 32'b01101110101001010000011111100011;
		#400 //0.31139365 * 1.21936884e-29 = 2.553728e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110111101110001111101111000;
		b = 32'b00000100010011100111010001100001;
		correct = 32'b01100010000110010011011011001000;
		#400 //1.7147598e-15 * 2.4268622e-36 = 7.065748e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010010001001110100010111100;
		b = 32'b11010000010011010001101101000101;
		correct = 32'b10100001011101011100010011000000;
		#400 //1.1461619e-08 * -13764466000.0 = -8.3269625e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101001010111111001101010010;
		b = 32'b01001011111011000001000100001001;
		correct = 32'b01000000101110100111100001010000;
		#400 //180303140.0 * 30941714.0 = 5.8271866
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100100100101101000010111000;
		b = 32'b11010110010111101000001000010111;
		correct = 32'b01010101101010001110100111110100;
		#400 //-1.4199105e+27 * -61162580000000.0 = 23215347000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111110000101001000000001011;
		b = 32'b01101110100010110010100011100110;
		correct = 32'b10100000101100101111010110111110;
		#400 //-6528440000.0 * 2.153393e+28 = -3.0316991e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110000111101110011010101110;
		b = 32'b01011111110011001001100001100100;
		correct = 32'b10110101110001101101001100111011;
		#400 //-43678400000000.0 * 2.9485287e+19 = -1.4813626e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000100111110001001110100001;
		b = 32'b10011101100101100001000011100001;
		correct = 32'b01101010100001111010111110010000;
		#400 //-325789.03 * -3.972212e-21 = 8.201703e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100010001100001110110101111;
		b = 32'b00010111111011011000110100110101;
		correct = 32'b01110011110101011000000001110100;
		#400 //51934908.0 * 1.5351412e-24 = 3.3830706e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011010001011011011111000110;
		b = 32'b11010010111100111100111100010001;
		correct = 32'b11001111110011111001101010110101;
		#400 //3.6472509e+21 * -523575530000.0 = -6966045000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011011010001011110100111101;
		b = 32'b01110001010100110110111011011000;
		correct = 32'b10100001100011001110011000001101;
		#400 //-999607300000.0 * 1.0469654e+30 = -9.547663e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100010100110011000001011101;
		b = 32'b10100010010111000011000010010110;
		correct = 32'b00111001011101011000100100001001;
		#400 //-6.987655e-22 * -2.984128e-18 = 0.0002341607
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010101101100001110000000100;
		b = 32'b01101010000000111111101101010001;
		correct = 32'b01000000001100001001110110001110;
		#400 //1.100784e+26 * 3.9889023e+25 = 2.7596164
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100101001010111101011111110;
		b = 32'b00110001001001101011110110001011;
		correct = 32'b01001010111111100001000011001000;
		#400 //0.020200249 * 2.4263922e-09 = 8325220.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101001101011010111110111010;
		b = 32'b00100100000110001100111111001111;
		correct = 32'b01101000100110000010111110110101;
		#400 //190512030.0 * 3.3135767e-17 = 5.749438e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110100110001101111111011111;
		b = 32'b10000111001111010100110010100100;
		correct = 32'b01001110110011101011110110011001;
		#400 //-2.4698207e-25 * -1.4241302e-34 = 1734266000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111110010100101111010001001;
		b = 32'b00000100011001100100101000111010;
		correct = 32'b11100010111000001111011001010011;
		#400 //-5.616876e-15 * 2.7070453e-36 = -2.0749101e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001011011111000110110100101;
		b = 32'b01000010110101100100001101000100;
		correct = 32'b01010110000011110001101111000111;
		#400 //4214266200000000.0 * 107.13138 = 39337366000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100000100111110110101111001;
		b = 32'b11010100110010001100110011010101;
		correct = 32'b00100110101111001001011111000111;
		#400 //-0.009028786 * -6899440000000.0 = 1.308626e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000111010111001111001101100;
		b = 32'b01101000101111011100100110010110;
		correct = 32'b11000111100111101110100100010100;
		#400 //-5.8336398e+29 * 7.169967e+24 = -81362.16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000001111101100000001101001;
		b = 32'b10000000111011111110110011101010;
		correct = 32'b01010110110010111000100000010111;
		#400 //-2.4654067e-24 * -2.2033672e-38 = 111892680000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110001000000001101100011110;
		b = 32'b00111011010000100111001101001111;
		correct = 32'b01000010010100101100100011001111;
		#400 //0.15635344 * 0.002967078 = 52.696102
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000110001011000101001100110011;
		b = 32'b10001111010011110010010111011000;
		correct = 32'b00110110010101001111011011111110;
		#400 //-3.241073e-35 * -1.02131764e-29 = 3.173423e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110000001001011001011000111;
		b = 32'b01110100011100000011000010111110;
		correct = 32'b00111001000011010110111011000110;
		#400 //1.0267037e+28 * 7.6119376e+31 = 0.00013488074
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100101110100010011001001110;
		b = 32'b00011110000100000001110100010001;
		correct = 32'b11011110001001010101011000000010;
		#400 //-0.022723343 * 7.629307e-21 = -2.978428e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001100110010100100001000010;
		b = 32'b01101000111100111001001000010110;
		correct = 32'b01010000001000010001101010101110;
		#400 //9.948587e+34 * 9.201839e+24 = 10811521000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101101100001010011101010011;
		b = 32'b01100001110011111101010111111011;
		correct = 32'b10010011010110011001011101101111;
		#400 //-1.316172e-06 * 4.7923687e+20 = -2.7463913e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101110000001111011001001010;
		b = 32'b10110110001111010111010111000000;
		correct = 32'b01001111000000100101110110110101;
		#400 //-6174.786 * -2.8231734e-06 = 2187179300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111110110010111100101101000;
		b = 32'b00101010101010100101010111111011;
		correct = 32'b01110100101000110110110000100101;
		#400 //3.1341341e+19 * 3.0257727e-13 = 1.0358128e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110111001001111010011110010000;
		b = 32'b01000110010001111100100101101001;
		correct = 32'b11110000010101101101001110101101;
		#400 //-3.400438e+33 * 12786.353 = -2.6594277e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100000011101000100110101111;
		b = 32'b00111110111100100010110000100001;
		correct = 32'b01000100100101101010110100101110;
		#400 //570.1513 * 0.47299293 = 1205.4119
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100100010111110100100101000;
		b = 32'b10110011111010100000011101000111;
		correct = 32'b11100000000110010000101111010010;
		#400 //4807297300000.0 * -1.0897798e-07 = -4.4112556e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101001000101100001001001010;
		b = 32'b11001110110111001111001101110110;
		correct = 32'b10110101101111001001001110111001;
		#400 //2604.143 * -1853471500.0 = -1.4050084e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011100000001100100110100000;
		b = 32'b01110110110110001000010110000111;
		correct = 32'b00111100000110000100010011111011;
		#400 //2.040721e+31 * 2.1957898e+33 = 0.00929379
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100011001001111011111100010;
		b = 32'b11000000000110110100011110001100;
		correct = 32'b01110011101111001011111001000000;
		#400 //-7.256295e+31 * -2.4262419 = 2.9907548e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101000000100001110100110110;
		b = 32'b01010011110001101110000011100110;
		correct = 32'b01000000101001110111110000110111;
		#400 //8941373000000.0 * 1708353400000.0 = 5.233913
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011011110000000010000110001;
		b = 32'b10100111111001100111000110101010;
		correct = 32'b00101011000010011100001010110100;
		#400 //-3.1304067e-27 * -6.396106e-15 = 4.894238e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100101001100010000110100111;
		b = 32'b11101001000100100101001001010010;
		correct = 32'b10001011000100010101010001010100;
		#400 //3.0944395e-07 * -1.1055745e+25 = -2.7989426e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101010001101001100100101010;
		b = 32'b00110000000010000010011001010110;
		correct = 32'b11101100101110101011010111100001;
		#400 //-8.944072e+17 * 4.953099e-10 = -1.8057528e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001101101001001010100001001;
		b = 32'b00110101000100011010011100101010;
		correct = 32'b01101100000111101011001000100000;
		#400 //4.1639413e+20 * 5.4259965e-07 = 7.674058e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111001101000111101101000000;
		b = 32'b01101000011000000001000000010101;
		correct = 32'b01010110010011100011010011101001;
		#400 //2.3990099e+38 * 4.232427e+24 = 56681660000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011011001010101000000100110;
		b = 32'b01001010010101000001000000100100;
		correct = 32'b10001000100010100110100101111010;
		#400 //-2.894338e-27 * 3474441.0 = -8.33037e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000110110101001010100110000;
		b = 32'b10100010001110111111100001101001;
		correct = 32'b11110110000101001101100010000101;
		#400 //1922674300000000.0 * -2.5474733e-18 = -7.547378e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111110100011111100010011001;
		b = 32'b10011100010100000101100101111011;
		correct = 32'b01101011000000001111111100000111;
		#400 //-107505.195 * -6.893708e-22 = 1.5594684e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010010011010011111110111001;
		b = 32'b11110011010110011101011111101101;
		correct = 32'b11000110011100010011001100001111;
		#400 //2.6642833e+35 * -1.7259337e+31 = -15436.765
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001100111011001110001011000;
		b = 32'b00001011101000111101100111001000;
		correct = 32'b11110101011101100100000000101011;
		#400 //-19.70134 * 6.3112997e-32 = -3.121598e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110000000111010100110011001;
		b = 32'b01100011000010010101011110010110;
		correct = 32'b11000010011101010110100111010100;
		#400 //-1.5543963e+23 * 2.5335152e+21 = -61.353348
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111010011110100010111110100;
		b = 32'b11110000100010110100111000010001;
		correct = 32'b00111110001111100111001111011000;
		#400 //-6.4147965e+28 * -3.4490234e+29 = 0.18598878
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101110001101001100100011100;
		b = 32'b10101110110011110001001111011001;
		correct = 32'b11110110011101011000010001101100;
		#400 //1.1723162e+23 * -9.416796e-11 = -1.2449205e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011010001101111000001001100;
		b = 32'b10001010110110110011010111101101;
		correct = 32'b11110111111010000101001101101010;
		#400 //198.93866 * -2.1109218e-32 = -9.4242555e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001101110111100001000001100010;
		b = 32'b10110110010000101001000101001110;
		correct = 32'b00010111000100100001011011001011;
		#400 //-1.368575e-30 * -2.8992831e-06 = 4.7203913e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010010001111001000100111100;
		b = 32'b00111100111111000100000101100100;
		correct = 32'b01101100110010101000011110011111;
		#400 //6.031552e+25 * 0.0307929 = 1.9587477e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101010100100110111111010100;
		b = 32'b11010101100111100011111001100111;
		correct = 32'b00111111001010100011011111000110;
		#400 //-14461109000000.0 * -21748857000000.0 = 0.66491354
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101010001111001010011010011;
		b = 32'b00010100010100010100100110000101;
		correct = 32'b11010000011101000010000010111001;
		#400 //-1.7310922e-16 * 1.0566303e-26 = -16383141000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100011011110100000110010100;
		b = 32'b10111101011100000111010010001000;
		correct = 32'b11010110011111101011100100110100;
		#400 //4110389600000.0 * -0.058704883 = -70017850000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101100110000100000011010011;
		b = 32'b01111010011010101001101010100011;
		correct = 32'b10100010101001100010001110000101;
		#400 //-1.3713751e+18 * 3.0453347e+35 = -4.5031998e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100111101110101010111110010;
		b = 32'b01001001100011001011000010110011;
		correct = 32'b10111010111000010000011010101110;
		#400 //-1978.6858 * 1152534.4 = -0.0017168128
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100000101110001011101011000;
		b = 32'b01100101110010100010010000010110;
		correct = 32'b00111101101111110101100100101111;
		#400 //1.1148562e+22 * 1.1932296e+23 = 0.09343182
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		$display ("Done.");
		$finish;
	end

endmodule
